netcdf ugrid-13x26x10-surface-subsurface-th-noice-dec-NGEE_SiteB.clm2.h0.0001-01-02-00000 {
dimensions:
	lndgrid = 338 ;
	gridcell = 338 ;
	landunit = 1352 ;
	column = 5408 ;
	pft = 10816 ;
	levgrnd = 15 ;
	levurb = 5 ;
	levlak = 10 ;
	numrad = 2 ;
	levsno = 5 ;
	ltype = 9 ;
	natpft = 17 ;
	string_length = 8 ;
	levdcmp = 15 ;
	hist_interval = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	float levlak(levlak) ;
		levlak:long_name = "coordinate lake levels" ;
		levlak:units = "m" ;
	float levdcmp(levdcmp) ;
		levdcmp:long_name = "coordinate soil levels" ;
		levdcmp:units = "m" ;
	float time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bounds" ;
	int mcdate(time) ;
		mcdate:long_name = "current date (YYYYMMDD)" ;
	int mcsec(time) ;
		mcsec:long_name = "current seconds of current date" ;
		mcsec:units = "s" ;
	int mdcur(time) ;
		mdcur:long_name = "current day (from base day)" ;
	int mscur(time) ;
		mscur:long_name = "current seconds of current day" ;
	int nstep(time) ;
		nstep:long_name = "time step" ;
	double time_bounds(time, hist_interval) ;
		time_bounds:long_name = "history time interval endpoints" ;
	char date_written(time, string_length) ;
	char time_written(time, string_length) ;
	float lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 1.e+36f ;
		lon:missing_value = 1.e+36f ;
	float lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 1.e+36f ;
		lat:missing_value = 1.e+36f ;
	float area(lndgrid) ;
		area:long_name = "grid cell areas" ;
		area:units = "km^2" ;
		area:_FillValue = 1.e+36f ;
		area:missing_value = 1.e+36f ;
	float topo(lndgrid) ;
		topo:long_name = "grid cell topography" ;
		topo:units = "m" ;
		topo:_FillValue = 1.e+36f ;
		topo:missing_value = 1.e+36f ;
	float landfrac(lndgrid) ;
		landfrac:long_name = "land fraction" ;
		landfrac:_FillValue = 1.e+36f ;
		landfrac:missing_value = 1.e+36f ;
	int landmask(lndgrid) ;
		landmask:long_name = "land/ocean mask (0.=ocean and 1.=land)" ;
		landmask:_FillValue = -9999 ;
		landmask:missing_value = -9999 ;
	int pftmask(lndgrid) ;
		pftmask:long_name = "pft real/fake mask (0.=fake and 1.=real)" ;
		pftmask:_FillValue = -9999 ;
		pftmask:missing_value = -9999 ;
	float ACTUAL_IMMOB(time, lndgrid) ;
		ACTUAL_IMMOB:long_name = "actual N immobilization" ;
		ACTUAL_IMMOB:units = "gN/m^2/s" ;
		ACTUAL_IMMOB:cell_methods = "time: mean" ;
		ACTUAL_IMMOB:_FillValue = 1.e+36f ;
		ACTUAL_IMMOB:missing_value = 1.e+36f ;
	float AGNPP(time, lndgrid) ;
		AGNPP:long_name = "aboveground NPP" ;
		AGNPP:units = "gC/m^2/s" ;
		AGNPP:cell_methods = "time: mean" ;
		AGNPP:_FillValue = 1.e+36f ;
		AGNPP:missing_value = 1.e+36f ;
	float ALT(time, lndgrid) ;
		ALT:long_name = "current active layer thickness" ;
		ALT:units = "m" ;
		ALT:cell_methods = "time: mean" ;
		ALT:_FillValue = 1.e+36f ;
		ALT:missing_value = 1.e+36f ;
	float ALTMAX(time, lndgrid) ;
		ALTMAX:long_name = "maximum annual active layer thickness" ;
		ALTMAX:units = "m" ;
		ALTMAX:cell_methods = "time: mean" ;
		ALTMAX:_FillValue = 1.e+36f ;
		ALTMAX:missing_value = 1.e+36f ;
	float ALTMAX_LASTYEAR(time, lndgrid) ;
		ALTMAX_LASTYEAR:long_name = "maximum prior year active layer thickness" ;
		ALTMAX_LASTYEAR:units = "m" ;
		ALTMAX_LASTYEAR:cell_methods = "time: mean" ;
		ALTMAX_LASTYEAR:_FillValue = 1.e+36f ;
		ALTMAX_LASTYEAR:missing_value = 1.e+36f ;
	float AR(time, lndgrid) ;
		AR:long_name = "autotrophic respiration (MR + GR)" ;
		AR:units = "gC/m^2/s" ;
		AR:cell_methods = "time: mean" ;
		AR:_FillValue = 1.e+36f ;
		AR:missing_value = 1.e+36f ;
	float BAF_CROP(time, lndgrid) ;
		BAF_CROP:long_name = "fractional area burned for crop" ;
		BAF_CROP:units = "proportion/sec" ;
		BAF_CROP:cell_methods = "time: mean" ;
		BAF_CROP:_FillValue = 1.e+36f ;
		BAF_CROP:missing_value = 1.e+36f ;
	float BAF_PEATF(time, lndgrid) ;
		BAF_PEATF:long_name = "fractional area burned in peatland" ;
		BAF_PEATF:units = "proportion/sec" ;
		BAF_PEATF:cell_methods = "time: mean" ;
		BAF_PEATF:_FillValue = 1.e+36f ;
		BAF_PEATF:missing_value = 1.e+36f ;
	float BCDEP(time, lndgrid) ;
		BCDEP:long_name = "total BC deposition (dry+wet) from atmosphere" ;
		BCDEP:units = "kg/m^2/s" ;
		BCDEP:cell_methods = "time: mean" ;
		BCDEP:_FillValue = 1.e+36f ;
		BCDEP:missing_value = 1.e+36f ;
	float BGNPP(time, lndgrid) ;
		BGNPP:long_name = "belowground NPP" ;
		BGNPP:units = "gC/m^2/s" ;
		BGNPP:cell_methods = "time: mean" ;
		BGNPP:_FillValue = 1.e+36f ;
		BGNPP:missing_value = 1.e+36f ;
	float BTRAN(time, lndgrid) ;
		BTRAN:long_name = "transpiration beta factor" ;
		BTRAN:units = "unitless" ;
		BTRAN:cell_methods = "time: mean" ;
		BTRAN:_FillValue = 1.e+36f ;
		BTRAN:missing_value = 1.e+36f ;
	float BUILDHEAT(time, lndgrid) ;
		BUILDHEAT:long_name = "heat flux from urban building interior to walls and roof" ;
		BUILDHEAT:units = "W/m^2" ;
		BUILDHEAT:cell_methods = "time: mean" ;
		BUILDHEAT:_FillValue = 1.e+36f ;
		BUILDHEAT:missing_value = 1.e+36f ;
	float CH4PROD(time, lndgrid) ;
		CH4PROD:long_name = "Gridcell total production of CH4" ;
		CH4PROD:units = "gC/m2/s" ;
		CH4PROD:cell_methods = "time: mean" ;
		CH4PROD:_FillValue = 1.e+36f ;
		CH4PROD:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_SAT(time, lndgrid) ;
		CH4_SURF_AERE_SAT:long_name = "aerenchyma surface CH4 flux for inundated area; (+ to atm)" ;
		CH4_SURF_AERE_SAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_SAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_UNSAT(time, lndgrid) ;
		CH4_SURF_AERE_UNSAT:long_name = "aerenchyma surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_AERE_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_SAT(time, lndgrid) ;
		CH4_SURF_DIFF_SAT:long_name = "diffusive surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_DIFF_SAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_SAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_UNSAT(time, lndgrid) ;
		CH4_SURF_DIFF_UNSAT:long_name = "diffusive surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_DIFF_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_SAT(time, lndgrid) ;
		CH4_SURF_EBUL_SAT:long_name = "ebullition surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_EBUL_SAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_SAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_UNSAT(time, lndgrid) ;
		CH4_SURF_EBUL_UNSAT:long_name = "ebullition surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_EBUL_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_UNSAT:missing_value = 1.e+36f ;
	float COL_CTRUNC(time, lndgrid) ;
		COL_CTRUNC:long_name = "column-level sink for C truncation" ;
		COL_CTRUNC:units = "gC/m^2" ;
		COL_CTRUNC:cell_methods = "time: mean" ;
		COL_CTRUNC:_FillValue = 1.e+36f ;
		COL_CTRUNC:missing_value = 1.e+36f ;
	float COL_FIRE_CLOSS(time, lndgrid) ;
		COL_FIRE_CLOSS:long_name = "total column-level fire C loss for non-peat fires outside land-type converted region" ;
		COL_FIRE_CLOSS:units = "gC/m^2/s" ;
		COL_FIRE_CLOSS:cell_methods = "time: mean" ;
		COL_FIRE_CLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_CLOSS:missing_value = 1.e+36f ;
	float COL_FIRE_NLOSS(time, lndgrid) ;
		COL_FIRE_NLOSS:long_name = "total column-level fire N loss" ;
		COL_FIRE_NLOSS:units = "gN/m^2/s" ;
		COL_FIRE_NLOSS:cell_methods = "time: mean" ;
		COL_FIRE_NLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_NLOSS:missing_value = 1.e+36f ;
	float COL_NTRUNC(time, lndgrid) ;
		COL_NTRUNC:long_name = "column-level sink for N truncation" ;
		COL_NTRUNC:units = "gN/m^2" ;
		COL_NTRUNC:cell_methods = "time: mean" ;
		COL_NTRUNC:_FillValue = 1.e+36f ;
		COL_NTRUNC:missing_value = 1.e+36f ;
	float CONC_CH4_SAT(time, levgrnd, lndgrid) ;
		CONC_CH4_SAT:long_name = "CH4 soil Concentration for inundated / lake area" ;
		CONC_CH4_SAT:units = "mol/m3" ;
		CONC_CH4_SAT:cell_methods = "time: mean" ;
		CONC_CH4_SAT:_FillValue = 1.e+36f ;
		CONC_CH4_SAT:missing_value = 1.e+36f ;
	float CONC_CH4_UNSAT(time, levgrnd, lndgrid) ;
		CONC_CH4_UNSAT:long_name = "CH4 soil Concentration for non-inundated area" ;
		CONC_CH4_UNSAT:units = "mol/m3" ;
		CONC_CH4_UNSAT:cell_methods = "time: mean" ;
		CONC_CH4_UNSAT:_FillValue = 1.e+36f ;
		CONC_CH4_UNSAT:missing_value = 1.e+36f ;
	float CONC_O2_SAT(time, levgrnd, lndgrid) ;
		CONC_O2_SAT:long_name = "O2 soil Concentration for inundated / lake area" ;
		CONC_O2_SAT:units = "mol/m3" ;
		CONC_O2_SAT:cell_methods = "time: mean" ;
		CONC_O2_SAT:_FillValue = 1.e+36f ;
		CONC_O2_SAT:missing_value = 1.e+36f ;
	float CONC_O2_UNSAT(time, levgrnd, lndgrid) ;
		CONC_O2_UNSAT:long_name = "O2 soil Concentration for non-inundated area" ;
		CONC_O2_UNSAT:units = "mol/m3" ;
		CONC_O2_UNSAT:cell_methods = "time: mean" ;
		CONC_O2_UNSAT:_FillValue = 1.e+36f ;
		CONC_O2_UNSAT:missing_value = 1.e+36f ;
	float CPOOL(time, lndgrid) ;
		CPOOL:long_name = "temporary photosynthate C pool" ;
		CPOOL:units = "gC/m^2" ;
		CPOOL:cell_methods = "time: mean" ;
		CPOOL:_FillValue = 1.e+36f ;
		CPOOL:missing_value = 1.e+36f ;
	float CWDC(time, lndgrid) ;
		CWDC:long_name = "CWD C" ;
		CWDC:units = "gC/m^2" ;
		CWDC:cell_methods = "time: mean" ;
		CWDC:_FillValue = 1.e+36f ;
		CWDC:missing_value = 1.e+36f ;
	float CWDC_HR(time, lndgrid) ;
		CWDC_HR:long_name = "coarse woody debris C heterotrophic respiration" ;
		CWDC_HR:units = "gC/m^2/s" ;
		CWDC_HR:cell_methods = "time: mean" ;
		CWDC_HR:_FillValue = 1.e+36f ;
		CWDC_HR:missing_value = 1.e+36f ;
	float CWDC_LOSS(time, lndgrid) ;
		CWDC_LOSS:long_name = "coarse woody debris C loss" ;
		CWDC_LOSS:units = "gC/m^2/s" ;
		CWDC_LOSS:cell_methods = "time: mean" ;
		CWDC_LOSS:_FillValue = 1.e+36f ;
		CWDC_LOSS:missing_value = 1.e+36f ;
	float CWDC_TO_LITR2C(time, lndgrid) ;
		CWDC_TO_LITR2C:long_name = "decomp. of coarse woody debris C to litter 2 C" ;
		CWDC_TO_LITR2C:units = "gC/m^2/s" ;
		CWDC_TO_LITR2C:cell_methods = "time: mean" ;
		CWDC_TO_LITR2C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR2C:missing_value = 1.e+36f ;
	float CWDC_TO_LITR3C(time, lndgrid) ;
		CWDC_TO_LITR3C:long_name = "decomp. of coarse woody debris C to litter 3 C" ;
		CWDC_TO_LITR3C:units = "gC/m^2/s" ;
		CWDC_TO_LITR3C:cell_methods = "time: mean" ;
		CWDC_TO_LITR3C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR3C:missing_value = 1.e+36f ;
	float CWDC_vr(time, levdcmp, lndgrid) ;
		CWDC_vr:long_name = "CWD C (vertically resolved)" ;
		CWDC_vr:units = "gC/m^3" ;
		CWDC_vr:cell_methods = "time: mean" ;
		CWDC_vr:_FillValue = 1.e+36f ;
		CWDC_vr:missing_value = 1.e+36f ;
	float CWDN(time, lndgrid) ;
		CWDN:long_name = "CWD N" ;
		CWDN:units = "gN/m^2" ;
		CWDN:cell_methods = "time: mean" ;
		CWDN:_FillValue = 1.e+36f ;
		CWDN:missing_value = 1.e+36f ;
	float CWDN_TO_LITR2N(time, lndgrid) ;
		CWDN_TO_LITR2N:long_name = "decomp. of coarse woody debris N to litter 2 N" ;
		CWDN_TO_LITR2N:units = "gN/m^2" ;
		CWDN_TO_LITR2N:cell_methods = "time: mean" ;
		CWDN_TO_LITR2N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR2N:missing_value = 1.e+36f ;
	float CWDN_TO_LITR3N(time, lndgrid) ;
		CWDN_TO_LITR3N:long_name = "decomp. of coarse woody debris N to litter 3 N" ;
		CWDN_TO_LITR3N:units = "gN/m^2" ;
		CWDN_TO_LITR3N:cell_methods = "time: mean" ;
		CWDN_TO_LITR3N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR3N:missing_value = 1.e+36f ;
	float CWDN_vr(time, levdcmp, lndgrid) ;
		CWDN_vr:long_name = "CWD N (vertically resolved)" ;
		CWDN_vr:units = "gN/m^3" ;
		CWDN_vr:cell_methods = "time: mean" ;
		CWDN_vr:_FillValue = 1.e+36f ;
		CWDN_vr:missing_value = 1.e+36f ;
	float DEADCROOTC(time, lndgrid) ;
		DEADCROOTC:long_name = "dead coarse root C" ;
		DEADCROOTC:units = "gC/m^2" ;
		DEADCROOTC:cell_methods = "time: mean" ;
		DEADCROOTC:_FillValue = 1.e+36f ;
		DEADCROOTC:missing_value = 1.e+36f ;
	float DEADCROOTN(time, lndgrid) ;
		DEADCROOTN:long_name = "dead coarse root N" ;
		DEADCROOTN:units = "gN/m^2" ;
		DEADCROOTN:cell_methods = "time: mean" ;
		DEADCROOTN:_FillValue = 1.e+36f ;
		DEADCROOTN:missing_value = 1.e+36f ;
	float DEADSTEMC(time, lndgrid) ;
		DEADSTEMC:long_name = "dead stem C" ;
		DEADSTEMC:units = "gC/m^2" ;
		DEADSTEMC:cell_methods = "time: mean" ;
		DEADSTEMC:_FillValue = 1.e+36f ;
		DEADSTEMC:missing_value = 1.e+36f ;
	float DEADSTEMN(time, lndgrid) ;
		DEADSTEMN:long_name = "dead stem N" ;
		DEADSTEMN:units = "gN/m^2" ;
		DEADSTEMN:cell_methods = "time: mean" ;
		DEADSTEMN:_FillValue = 1.e+36f ;
		DEADSTEMN:missing_value = 1.e+36f ;
	float DENIT(time, lndgrid) ;
		DENIT:long_name = "total rate of denitrification" ;
		DENIT:units = "gN/m^2/s" ;
		DENIT:cell_methods = "time: mean" ;
		DENIT:_FillValue = 1.e+36f ;
		DENIT:missing_value = 1.e+36f ;
	float DISPVEGC(time, lndgrid) ;
		DISPVEGC:long_name = "displayed veg carbon, excluding storage and cpool" ;
		DISPVEGC:units = "gC/m^2" ;
		DISPVEGC:cell_methods = "time: mean" ;
		DISPVEGC:_FillValue = 1.e+36f ;
		DISPVEGC:missing_value = 1.e+36f ;
	float DISPVEGN(time, lndgrid) ;
		DISPVEGN:long_name = "displayed vegetation nitrogen" ;
		DISPVEGN:units = "gN/m^2" ;
		DISPVEGN:cell_methods = "time: mean" ;
		DISPVEGN:_FillValue = 1.e+36f ;
		DISPVEGN:missing_value = 1.e+36f ;
	float DSTDEP(time, lndgrid) ;
		DSTDEP:long_name = "total dust deposition (dry+wet) from atmosphere" ;
		DSTDEP:units = "kg/m^2/s" ;
		DSTDEP:cell_methods = "time: mean" ;
		DSTDEP:_FillValue = 1.e+36f ;
		DSTDEP:missing_value = 1.e+36f ;
	float DSTFLXT(time, lndgrid) ;
		DSTFLXT:long_name = "total surface dust emission" ;
		DSTFLXT:units = "kg/m2/s" ;
		DSTFLXT:cell_methods = "time: mean" ;
		DSTFLXT:_FillValue = 1.e+36f ;
		DSTFLXT:missing_value = 1.e+36f ;
	float DWT_CLOSS(time, lndgrid) ;
		DWT_CLOSS:long_name = "total carbon loss from land cover conversion" ;
		DWT_CLOSS:units = "gC/m^2/s" ;
		DWT_CLOSS:cell_methods = "time: mean" ;
		DWT_CLOSS:_FillValue = 1.e+36f ;
		DWT_CLOSS:missing_value = 1.e+36f ;
	float DWT_CONV_CFLUX(time, lndgrid) ;
		DWT_CONV_CFLUX:long_name = "conversion C flux (immediate loss to atm)" ;
		DWT_CONV_CFLUX:units = "gC/m^2/s" ;
		DWT_CONV_CFLUX:cell_methods = "time: mean" ;
		DWT_CONV_CFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_CFLUX:missing_value = 1.e+36f ;
	float DWT_CONV_NFLUX(time, lndgrid) ;
		DWT_CONV_NFLUX:long_name = "conversion N flux (immediate loss to atm)" ;
		DWT_CONV_NFLUX:units = "gN/m^2/s" ;
		DWT_CONV_NFLUX:cell_methods = "time: mean" ;
		DWT_CONV_NFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_NFLUX:missing_value = 1.e+36f ;
	float DWT_NLOSS(time, lndgrid) ;
		DWT_NLOSS:long_name = "total nitrogen loss from landcover conversion" ;
		DWT_NLOSS:units = "gN/m^2/s" ;
		DWT_NLOSS:cell_methods = "time: mean" ;
		DWT_NLOSS:_FillValue = 1.e+36f ;
		DWT_NLOSS:missing_value = 1.e+36f ;
	float DWT_PROD100C_GAIN(time, lndgrid) ;
		DWT_PROD100C_GAIN:long_name = "landcover change-driven addition to 100-yr wood product pool" ;
		DWT_PROD100C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD100C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD100N_GAIN(time, lndgrid) ;
		DWT_PROD100N_GAIN:long_name = "addition to 100-yr wood product pool" ;
		DWT_PROD100N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD100N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100N_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10C_GAIN(time, lndgrid) ;
		DWT_PROD10C_GAIN:long_name = "landcover change-driven addition to 10-yr wood product pool" ;
		DWT_PROD10C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD10C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10N_GAIN(time, lndgrid) ;
		DWT_PROD10N_GAIN:long_name = "addition to 10-yr wood product pool" ;
		DWT_PROD10N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD10N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10N_GAIN:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDC_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDC_TO_DEADSTEM:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_LEAF(time, lndgrid) ;
		DWT_SEEDC_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDC_TO_LEAF:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_LEAF:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDN_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDN_TO_DEADSTEM:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_LEAF(time, lndgrid) ;
		DWT_SEEDN_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDN_TO_LEAF:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_LEAF:missing_value = 1.e+36f ;
	float EFLX_DYNBAL(time, lndgrid) ;
		EFLX_DYNBAL:long_name = "dynamic land cover change conversion energy flux" ;
		EFLX_DYNBAL:units = "W/m^2" ;
		EFLX_DYNBAL:cell_methods = "time: mean" ;
		EFLX_DYNBAL:_FillValue = 1.e+36f ;
		EFLX_DYNBAL:missing_value = 1.e+36f ;
	float EFLX_GRND_LAKE(time, lndgrid) ;
		EFLX_GRND_LAKE:long_name = "net heat flux into lake/snow surface, excluding light transmission" ;
		EFLX_GRND_LAKE:units = "W/m^2" ;
		EFLX_GRND_LAKE:cell_methods = "time: mean" ;
		EFLX_GRND_LAKE:_FillValue = 1.e+36f ;
		EFLX_GRND_LAKE:missing_value = 1.e+36f ;
	float EFLX_LH_TOT(time, lndgrid) ;
		EFLX_LH_TOT:long_name = "total latent heat flux [+ to atm]" ;
		EFLX_LH_TOT:units = "W/m^2" ;
		EFLX_LH_TOT:cell_methods = "time: mean" ;
		EFLX_LH_TOT:_FillValue = 1.e+36f ;
		EFLX_LH_TOT:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_R(time, lndgrid) ;
		EFLX_LH_TOT_R:long_name = "Rural total evaporation" ;
		EFLX_LH_TOT_R:units = "W/m^2" ;
		EFLX_LH_TOT_R:cell_methods = "time: mean" ;
		EFLX_LH_TOT_R:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_R:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_U(time, lndgrid) ;
		EFLX_LH_TOT_U:long_name = "Urban total evaporation" ;
		EFLX_LH_TOT_U:units = "W/m^2" ;
		EFLX_LH_TOT_U:cell_methods = "time: mean" ;
		EFLX_LH_TOT_U:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_U:missing_value = 1.e+36f ;
	float ELAI(time, lndgrid) ;
		ELAI:long_name = "exposed one-sided leaf area index" ;
		ELAI:units = "m^2/m^2" ;
		ELAI:cell_methods = "time: mean" ;
		ELAI:_FillValue = 1.e+36f ;
		ELAI:missing_value = 1.e+36f ;
	float ER(time, lndgrid) ;
		ER:long_name = "total ecosystem respiration, autotrophic + heterotrophic" ;
		ER:units = "gC/m^2/s" ;
		ER:cell_methods = "time: mean" ;
		ER:_FillValue = 1.e+36f ;
		ER:missing_value = 1.e+36f ;
	float ERRH2O(time, lndgrid) ;
		ERRH2O:long_name = "total water conservation error" ;
		ERRH2O:units = "mm" ;
		ERRH2O:cell_methods = "time: mean" ;
		ERRH2O:_FillValue = 1.e+36f ;
		ERRH2O:missing_value = 1.e+36f ;
	float ERRH2OSNO(time, lndgrid) ;
		ERRH2OSNO:long_name = "imbalance in snow depth (liquid water)" ;
		ERRH2OSNO:units = "mm" ;
		ERRH2OSNO:cell_methods = "time: mean" ;
		ERRH2OSNO:_FillValue = 1.e+36f ;
		ERRH2OSNO:missing_value = 1.e+36f ;
	float ERRSEB(time, lndgrid) ;
		ERRSEB:long_name = "surface energy conservation error" ;
		ERRSEB:units = "W/m^2" ;
		ERRSEB:cell_methods = "time: mean" ;
		ERRSEB:_FillValue = 1.e+36f ;
		ERRSEB:missing_value = 1.e+36f ;
	float ERRSOI(time, lndgrid) ;
		ERRSOI:long_name = "soil/lake energy conservation error" ;
		ERRSOI:units = "W/m^2" ;
		ERRSOI:cell_methods = "time: mean" ;
		ERRSOI:_FillValue = 1.e+36f ;
		ERRSOI:missing_value = 1.e+36f ;
	float ERRSOL(time, lndgrid) ;
		ERRSOL:long_name = "solar radiation conservation error" ;
		ERRSOL:units = "W/m^2" ;
		ERRSOL:cell_methods = "time: mean" ;
		ERRSOL:_FillValue = 1.e+36f ;
		ERRSOL:missing_value = 1.e+36f ;
	float ESAI(time, lndgrid) ;
		ESAI:long_name = "exposed one-sided stem area index" ;
		ESAI:units = "m^2/m^2" ;
		ESAI:cell_methods = "time: mean" ;
		ESAI:_FillValue = 1.e+36f ;
		ESAI:missing_value = 1.e+36f ;
	float FAREA_BURNED(time, lndgrid) ;
		FAREA_BURNED:long_name = "fractional area burned" ;
		FAREA_BURNED:units = "proportion/sec" ;
		FAREA_BURNED:cell_methods = "time: mean" ;
		FAREA_BURNED:_FillValue = 1.e+36f ;
		FAREA_BURNED:missing_value = 1.e+36f ;
	float FCEV(time, lndgrid) ;
		FCEV:long_name = "canopy evaporation" ;
		FCEV:units = "W/m^2" ;
		FCEV:cell_methods = "time: mean" ;
		FCEV:_FillValue = 1.e+36f ;
		FCEV:missing_value = 1.e+36f ;
	float FCH4(time, lndgrid) ;
		FCH4:long_name = "Gridcell surface CH4 flux to atmosphere (+ to atm)" ;
		FCH4:units = "kgC/m2/s" ;
		FCH4:cell_methods = "time: mean" ;
		FCH4:_FillValue = 1.e+36f ;
		FCH4:missing_value = 1.e+36f ;
	float FCH4TOCO2(time, lndgrid) ;
		FCH4TOCO2:long_name = "Gridcell oxidation of CH4 to CO2" ;
		FCH4TOCO2:units = "gC/m2/s" ;
		FCH4TOCO2:cell_methods = "time: mean" ;
		FCH4TOCO2:_FillValue = 1.e+36f ;
		FCH4TOCO2:missing_value = 1.e+36f ;
	float FCH4_DFSAT(time, lndgrid) ;
		FCH4_DFSAT:long_name = "CH4 additional flux due to changing fsat, vegetated landunits only" ;
		FCH4_DFSAT:units = "kgC/m2/s" ;
		FCH4_DFSAT:cell_methods = "time: mean" ;
		FCH4_DFSAT:_FillValue = 1.e+36f ;
		FCH4_DFSAT:missing_value = 1.e+36f ;
	float FCOV(time, lndgrid) ;
		FCOV:long_name = "fractional impermeable area" ;
		FCOV:units = "unitless" ;
		FCOV:cell_methods = "time: mean" ;
		FCOV:_FillValue = 1.e+36f ;
		FCOV:missing_value = 1.e+36f ;
	float FCTR(time, lndgrid) ;
		FCTR:long_name = "canopy transpiration" ;
		FCTR:units = "W/m^2" ;
		FCTR:cell_methods = "time: mean" ;
		FCTR:_FillValue = 1.e+36f ;
		FCTR:missing_value = 1.e+36f ;
	float FGEV(time, lndgrid) ;
		FGEV:long_name = "ground evaporation" ;
		FGEV:units = "W/m^2" ;
		FGEV:cell_methods = "time: mean" ;
		FGEV:_FillValue = 1.e+36f ;
		FGEV:missing_value = 1.e+36f ;
	float FGR(time, lndgrid) ;
		FGR:long_name = "heat flux into soil/snow including snow melt and lake / snow light transmission" ;
		FGR:units = "W/m^2" ;
		FGR:cell_methods = "time: mean" ;
		FGR:_FillValue = 1.e+36f ;
		FGR:missing_value = 1.e+36f ;
	float FGR12(time, lndgrid) ;
		FGR12:long_name = "heat flux between soil layers 1 and 2" ;
		FGR12:units = "W/m^2" ;
		FGR12:cell_methods = "time: mean" ;
		FGR12:_FillValue = 1.e+36f ;
		FGR12:missing_value = 1.e+36f ;
	float FGR_R(time, lndgrid) ;
		FGR_R:long_name = "Rural heat flux into soil/snow including snow melt and snow light transmission" ;
		FGR_R:units = "W/m^2" ;
		FGR_R:cell_methods = "time: mean" ;
		FGR_R:_FillValue = 1.e+36f ;
		FGR_R:missing_value = 1.e+36f ;
	float FGR_U(time, lndgrid) ;
		FGR_U:long_name = "Urban heat flux into soil/snow including snow melt" ;
		FGR_U:units = "W/m^2" ;
		FGR_U:cell_methods = "time: mean" ;
		FGR_U:_FillValue = 1.e+36f ;
		FGR_U:missing_value = 1.e+36f ;
	float FH2OSFC(time, lndgrid) ;
		FH2OSFC:long_name = "fraction of ground covered by surface water" ;
		FH2OSFC:units = "unitless" ;
		FH2OSFC:cell_methods = "time: mean" ;
		FH2OSFC:_FillValue = 1.e+36f ;
		FH2OSFC:missing_value = 1.e+36f ;
	float FINUNDATED(time, lndgrid) ;
		FINUNDATED:long_name = "fractional inundated area of vegetated columns" ;
		FINUNDATED:units = "unitless" ;
		FINUNDATED:cell_methods = "time: mean" ;
		FINUNDATED:_FillValue = 1.e+36f ;
		FINUNDATED:missing_value = 1.e+36f ;
	float FINUNDATED_LAG(time, lndgrid) ;
		FINUNDATED_LAG:long_name = "time-lagged inundated fraction of vegetated columns" ;
		FINUNDATED_LAG:units = "unitless" ;
		FINUNDATED_LAG:cell_methods = "time: mean" ;
		FINUNDATED_LAG:_FillValue = 1.e+36f ;
		FINUNDATED_LAG:missing_value = 1.e+36f ;
	float FIRA(time, lndgrid) ;
		FIRA:long_name = "net infrared (longwave) radiation" ;
		FIRA:units = "W/m^2" ;
		FIRA:cell_methods = "time: mean" ;
		FIRA:_FillValue = 1.e+36f ;
		FIRA:missing_value = 1.e+36f ;
	float FIRA_R(time, lndgrid) ;
		FIRA_R:long_name = "Rural net infrared (longwave) radiation" ;
		FIRA_R:units = "W/m^2" ;
		FIRA_R:cell_methods = "time: mean" ;
		FIRA_R:_FillValue = 1.e+36f ;
		FIRA_R:missing_value = 1.e+36f ;
	float FIRA_U(time, lndgrid) ;
		FIRA_U:long_name = "Urban net infrared (longwave) radiation" ;
		FIRA_U:units = "W/m^2" ;
		FIRA_U:cell_methods = "time: mean" ;
		FIRA_U:_FillValue = 1.e+36f ;
		FIRA_U:missing_value = 1.e+36f ;
	float FIRE(time, lndgrid) ;
		FIRE:long_name = "emitted infrared (longwave) radiation" ;
		FIRE:units = "W/m^2" ;
		FIRE:cell_methods = "time: mean" ;
		FIRE:_FillValue = 1.e+36f ;
		FIRE:missing_value = 1.e+36f ;
	float FIRE_R(time, lndgrid) ;
		FIRE_R:long_name = "Rural emitted infrared (longwave) radiation" ;
		FIRE_R:units = "W/m^2" ;
		FIRE_R:cell_methods = "time: mean" ;
		FIRE_R:_FillValue = 1.e+36f ;
		FIRE_R:missing_value = 1.e+36f ;
	float FIRE_U(time, lndgrid) ;
		FIRE_U:long_name = "Urban emitted infrared (longwave) radiation" ;
		FIRE_U:units = "W/m^2" ;
		FIRE_U:cell_methods = "time: mean" ;
		FIRE_U:_FillValue = 1.e+36f ;
		FIRE_U:missing_value = 1.e+36f ;
	float FLDS(time, lndgrid) ;
		FLDS:long_name = "atmospheric longwave radiation" ;
		FLDS:units = "W/m^2" ;
		FLDS:cell_methods = "time: mean" ;
		FLDS:_FillValue = 1.e+36f ;
		FLDS:missing_value = 1.e+36f ;
	float FPG(time, lndgrid) ;
		FPG:long_name = "fraction of potential gpp" ;
		FPG:units = "proportion" ;
		FPG:cell_methods = "time: mean" ;
		FPG:_FillValue = 1.e+36f ;
		FPG:missing_value = 1.e+36f ;
	float FPI(time, lndgrid) ;
		FPI:long_name = "fraction of potential immobilization" ;
		FPI:units = "proportion" ;
		FPI:cell_methods = "time: mean" ;
		FPI:_FillValue = 1.e+36f ;
		FPI:missing_value = 1.e+36f ;
	float FPI_vr(time, levdcmp, lndgrid) ;
		FPI_vr:long_name = "fraction of potential immobilization" ;
		FPI_vr:units = "proportion" ;
		FPI_vr:cell_methods = "time: mean" ;
		FPI_vr:_FillValue = 1.e+36f ;
		FPI_vr:missing_value = 1.e+36f ;
	float FPSN(time, lndgrid) ;
		FPSN:long_name = "photosynthesis" ;
		FPSN:units = "umol/m2s" ;
		FPSN:cell_methods = "time: mean" ;
		FPSN:_FillValue = 1.e+36f ;
		FPSN:missing_value = 1.e+36f ;
	float FPSN_WC(time, lndgrid) ;
		FPSN_WC:long_name = "Rubisco-limited photosynthesis" ;
		FPSN_WC:units = "umol/m2s" ;
		FPSN_WC:cell_methods = "time: mean" ;
		FPSN_WC:_FillValue = 1.e+36f ;
		FPSN_WC:missing_value = 1.e+36f ;
	float FPSN_WJ(time, lndgrid) ;
		FPSN_WJ:long_name = "RuBP-limited photosynthesis" ;
		FPSN_WJ:units = "umol/m2s" ;
		FPSN_WJ:cell_methods = "time: mean" ;
		FPSN_WJ:_FillValue = 1.e+36f ;
		FPSN_WJ:missing_value = 1.e+36f ;
	float FPSN_WP(time, lndgrid) ;
		FPSN_WP:long_name = "Product-limited photosynthesis" ;
		FPSN_WP:units = "umol/m2s" ;
		FPSN_WP:cell_methods = "time: mean" ;
		FPSN_WP:_FillValue = 1.e+36f ;
		FPSN_WP:missing_value = 1.e+36f ;
	float FROOTC(time, lndgrid) ;
		FROOTC:long_name = "fine root C" ;
		FROOTC:units = "gC/m^2" ;
		FROOTC:cell_methods = "time: mean" ;
		FROOTC:_FillValue = 1.e+36f ;
		FROOTC:missing_value = 1.e+36f ;
	float FROOTC_ALLOC(time, lndgrid) ;
		FROOTC_ALLOC:long_name = "fine root C allocation" ;
		FROOTC_ALLOC:units = "gC/m^2/s" ;
		FROOTC_ALLOC:cell_methods = "time: mean" ;
		FROOTC_ALLOC:_FillValue = 1.e+36f ;
		FROOTC_ALLOC:missing_value = 1.e+36f ;
	float FROOTC_LOSS(time, lndgrid) ;
		FROOTC_LOSS:long_name = "fine root C loss" ;
		FROOTC_LOSS:units = "gC/m^2/s" ;
		FROOTC_LOSS:cell_methods = "time: mean" ;
		FROOTC_LOSS:_FillValue = 1.e+36f ;
		FROOTC_LOSS:missing_value = 1.e+36f ;
	float FROOTN(time, lndgrid) ;
		FROOTN:long_name = "fine root N" ;
		FROOTN:units = "gN/m^2" ;
		FROOTN:cell_methods = "time: mean" ;
		FROOTN:_FillValue = 1.e+36f ;
		FROOTN:missing_value = 1.e+36f ;
	float FROST_TABLE(time, lndgrid) ;
		FROST_TABLE:long_name = "frost table depth (vegetated landunits only)" ;
		FROST_TABLE:units = "m" ;
		FROST_TABLE:cell_methods = "time: mean" ;
		FROST_TABLE:_FillValue = 1.e+36f ;
		FROST_TABLE:missing_value = 1.e+36f ;
	float FSA(time, lndgrid) ;
		FSA:long_name = "absorbed solar radiation" ;
		FSA:units = "W/m^2" ;
		FSA:cell_methods = "time: mean" ;
		FSA:_FillValue = 1.e+36f ;
		FSA:missing_value = 1.e+36f ;
	float FSAT(time, lndgrid) ;
		FSAT:long_name = "fractional area with water table at surface" ;
		FSAT:units = "unitless" ;
		FSAT:cell_methods = "time: mean" ;
		FSAT:_FillValue = 1.e+36f ;
		FSAT:missing_value = 1.e+36f ;
	float FSA_R(time, lndgrid) ;
		FSA_R:long_name = "Rural absorbed solar radiation" ;
		FSA_R:units = "W/m^2" ;
		FSA_R:cell_methods = "time: mean" ;
		FSA_R:_FillValue = 1.e+36f ;
		FSA_R:missing_value = 1.e+36f ;
	float FSA_U(time, lndgrid) ;
		FSA_U:long_name = "Urban absorbed solar radiation" ;
		FSA_U:units = "W/m^2" ;
		FSA_U:cell_methods = "time: mean" ;
		FSA_U:_FillValue = 1.e+36f ;
		FSA_U:missing_value = 1.e+36f ;
	float FSDS(time, lndgrid) ;
		FSDS:long_name = "atmospheric incident solar radiation" ;
		FSDS:units = "W/m^2" ;
		FSDS:cell_methods = "time: mean" ;
		FSDS:_FillValue = 1.e+36f ;
		FSDS:missing_value = 1.e+36f ;
	float FSDSND(time, lndgrid) ;
		FSDSND:long_name = "direct nir incident solar radiation" ;
		FSDSND:units = "W/m^2" ;
		FSDSND:cell_methods = "time: mean" ;
		FSDSND:_FillValue = 1.e+36f ;
		FSDSND:missing_value = 1.e+36f ;
	float FSDSNDLN(time, lndgrid) ;
		FSDSNDLN:long_name = "direct nir incident solar radiation at local noon" ;
		FSDSNDLN:units = "W/m^2" ;
		FSDSNDLN:cell_methods = "time: mean" ;
		FSDSNDLN:_FillValue = 1.e+36f ;
		FSDSNDLN:missing_value = 1.e+36f ;
	float FSDSNI(time, lndgrid) ;
		FSDSNI:long_name = "diffuse nir incident solar radiation" ;
		FSDSNI:units = "W/m^2" ;
		FSDSNI:cell_methods = "time: mean" ;
		FSDSNI:_FillValue = 1.e+36f ;
		FSDSNI:missing_value = 1.e+36f ;
	float FSDSVD(time, lndgrid) ;
		FSDSVD:long_name = "direct vis incident solar radiation" ;
		FSDSVD:units = "W/m^2" ;
		FSDSVD:cell_methods = "time: mean" ;
		FSDSVD:_FillValue = 1.e+36f ;
		FSDSVD:missing_value = 1.e+36f ;
	float FSDSVDLN(time, lndgrid) ;
		FSDSVDLN:long_name = "direct vis incident solar radiation at local noon" ;
		FSDSVDLN:units = "W/m^2" ;
		FSDSVDLN:cell_methods = "time: mean" ;
		FSDSVDLN:_FillValue = 1.e+36f ;
		FSDSVDLN:missing_value = 1.e+36f ;
	float FSDSVI(time, lndgrid) ;
		FSDSVI:long_name = "diffuse vis incident solar radiation" ;
		FSDSVI:units = "W/m^2" ;
		FSDSVI:cell_methods = "time: mean" ;
		FSDSVI:_FillValue = 1.e+36f ;
		FSDSVI:missing_value = 1.e+36f ;
	float FSDSVILN(time, lndgrid) ;
		FSDSVILN:long_name = "diffuse vis incident solar radiation at local noon" ;
		FSDSVILN:units = "W/m^2" ;
		FSDSVILN:cell_methods = "time: mean" ;
		FSDSVILN:_FillValue = 1.e+36f ;
		FSDSVILN:missing_value = 1.e+36f ;
	float FSH(time, lndgrid) ;
		FSH:long_name = "sensible heat" ;
		FSH:units = "W/m^2" ;
		FSH:cell_methods = "time: mean" ;
		FSH:_FillValue = 1.e+36f ;
		FSH:missing_value = 1.e+36f ;
	float FSH_G(time, lndgrid) ;
		FSH_G:long_name = "sensible heat from ground" ;
		FSH_G:units = "W/m^2" ;
		FSH_G:cell_methods = "time: mean" ;
		FSH_G:_FillValue = 1.e+36f ;
		FSH_G:missing_value = 1.e+36f ;
	float FSH_NODYNLNDUSE(time, lndgrid) ;
		FSH_NODYNLNDUSE:long_name = "sensible heat not including correction for land use change" ;
		FSH_NODYNLNDUSE:units = "W/m^2" ;
		FSH_NODYNLNDUSE:cell_methods = "time: mean" ;
		FSH_NODYNLNDUSE:_FillValue = 1.e+36f ;
		FSH_NODYNLNDUSE:missing_value = 1.e+36f ;
	float FSH_R(time, lndgrid) ;
		FSH_R:long_name = "Rural sensible heat" ;
		FSH_R:units = "W/m^2" ;
		FSH_R:cell_methods = "time: mean" ;
		FSH_R:_FillValue = 1.e+36f ;
		FSH_R:missing_value = 1.e+36f ;
	float FSH_U(time, lndgrid) ;
		FSH_U:long_name = "Urban sensible heat" ;
		FSH_U:units = "W/m^2" ;
		FSH_U:cell_methods = "time: mean" ;
		FSH_U:_FillValue = 1.e+36f ;
		FSH_U:missing_value = 1.e+36f ;
	float FSH_V(time, lndgrid) ;
		FSH_V:long_name = "sensible heat from veg" ;
		FSH_V:units = "W/m^2" ;
		FSH_V:cell_methods = "time: mean" ;
		FSH_V:_FillValue = 1.e+36f ;
		FSH_V:missing_value = 1.e+36f ;
	float FSM(time, lndgrid) ;
		FSM:long_name = "snow melt heat flux" ;
		FSM:units = "W/m^2" ;
		FSM:cell_methods = "time: mean" ;
		FSM:_FillValue = 1.e+36f ;
		FSM:missing_value = 1.e+36f ;
	float FSM_R(time, lndgrid) ;
		FSM_R:long_name = "Rural snow melt heat flux" ;
		FSM_R:units = "W/m^2" ;
		FSM_R:cell_methods = "time: mean" ;
		FSM_R:_FillValue = 1.e+36f ;
		FSM_R:missing_value = 1.e+36f ;
	float FSM_U(time, lndgrid) ;
		FSM_U:long_name = "Urban snow melt heat flux" ;
		FSM_U:units = "W/m^2" ;
		FSM_U:cell_methods = "time: mean" ;
		FSM_U:_FillValue = 1.e+36f ;
		FSM_U:missing_value = 1.e+36f ;
	float FSNO(time, lndgrid) ;
		FSNO:long_name = "fraction of ground covered by snow" ;
		FSNO:units = "unitless" ;
		FSNO:cell_methods = "time: mean" ;
		FSNO:_FillValue = 1.e+36f ;
		FSNO:missing_value = 1.e+36f ;
	float FSNO_EFF(time, lndgrid) ;
		FSNO_EFF:long_name = "effective fraction of ground covered by snow" ;
		FSNO_EFF:units = "unitless" ;
		FSNO_EFF:cell_methods = "time: mean" ;
		FSNO_EFF:_FillValue = 1.e+36f ;
		FSNO_EFF:missing_value = 1.e+36f ;
	float FSR(time, lndgrid) ;
		FSR:long_name = "reflected solar radiation" ;
		FSR:units = "W/m^2" ;
		FSR:cell_methods = "time: mean" ;
		FSR:_FillValue = 1.e+36f ;
		FSR:missing_value = 1.e+36f ;
	float FSRND(time, lndgrid) ;
		FSRND:long_name = "direct nir reflected solar radiation" ;
		FSRND:units = "W/m^2" ;
		FSRND:cell_methods = "time: mean" ;
		FSRND:_FillValue = 1.e+36f ;
		FSRND:missing_value = 1.e+36f ;
	float FSRNDLN(time, lndgrid) ;
		FSRNDLN:long_name = "direct nir reflected solar radiation at local noon" ;
		FSRNDLN:units = "W/m^2" ;
		FSRNDLN:cell_methods = "time: mean" ;
		FSRNDLN:_FillValue = 1.e+36f ;
		FSRNDLN:missing_value = 1.e+36f ;
	float FSRNI(time, lndgrid) ;
		FSRNI:long_name = "diffuse nir reflected solar radiation" ;
		FSRNI:units = "W/m^2" ;
		FSRNI:cell_methods = "time: mean" ;
		FSRNI:_FillValue = 1.e+36f ;
		FSRNI:missing_value = 1.e+36f ;
	float FSRVD(time, lndgrid) ;
		FSRVD:long_name = "direct vis reflected solar radiation" ;
		FSRVD:units = "W/m^2" ;
		FSRVD:cell_methods = "time: mean" ;
		FSRVD:_FillValue = 1.e+36f ;
		FSRVD:missing_value = 1.e+36f ;
	float FSRVDLN(time, lndgrid) ;
		FSRVDLN:long_name = "direct vis reflected solar radiation at local noon" ;
		FSRVDLN:units = "W/m^2" ;
		FSRVDLN:cell_methods = "time: mean" ;
		FSRVDLN:_FillValue = 1.e+36f ;
		FSRVDLN:missing_value = 1.e+36f ;
	float FSRVI(time, lndgrid) ;
		FSRVI:long_name = "diffuse vis reflected solar radiation" ;
		FSRVI:units = "W/m^2" ;
		FSRVI:cell_methods = "time: mean" ;
		FSRVI:_FillValue = 1.e+36f ;
		FSRVI:missing_value = 1.e+36f ;
	float FUELC(time, lndgrid) ;
		FUELC:long_name = "fuel load" ;
		FUELC:units = "gC/m^2" ;
		FUELC:cell_methods = "time: mean" ;
		FUELC:_FillValue = 1.e+36f ;
		FUELC:missing_value = 1.e+36f ;
	float F_DENIT(time, lndgrid) ;
		F_DENIT:long_name = "denitrification flux" ;
		F_DENIT:units = "gN/m^2/s" ;
		F_DENIT:cell_methods = "time: mean" ;
		F_DENIT:_FillValue = 1.e+36f ;
		F_DENIT:missing_value = 1.e+36f ;
	float F_DENIT_vr(time, levdcmp, lndgrid) ;
		F_DENIT_vr:long_name = "denitrification flux" ;
		F_DENIT_vr:units = "gN/m^3/s" ;
		F_DENIT_vr:cell_methods = "time: mean" ;
		F_DENIT_vr:_FillValue = 1.e+36f ;
		F_DENIT_vr:missing_value = 1.e+36f ;
	float F_N2O_DENIT(time, lndgrid) ;
		F_N2O_DENIT:long_name = "denitrification N2O flux" ;
		F_N2O_DENIT:units = "gN/m^2/s" ;
		F_N2O_DENIT:cell_methods = "time: mean" ;
		F_N2O_DENIT:_FillValue = 1.e+36f ;
		F_N2O_DENIT:missing_value = 1.e+36f ;
	float F_N2O_NIT(time, lndgrid) ;
		F_N2O_NIT:long_name = "nitrification N2O flux" ;
		F_N2O_NIT:units = "gN/m^2/s" ;
		F_N2O_NIT:cell_methods = "time: mean" ;
		F_N2O_NIT:_FillValue = 1.e+36f ;
		F_N2O_NIT:missing_value = 1.e+36f ;
	float F_NIT(time, lndgrid) ;
		F_NIT:long_name = "nitrification flux" ;
		F_NIT:units = "gN/m^2/s" ;
		F_NIT:cell_methods = "time: mean" ;
		F_NIT:_FillValue = 1.e+36f ;
		F_NIT:missing_value = 1.e+36f ;
	float F_NIT_vr(time, levdcmp, lndgrid) ;
		F_NIT_vr:long_name = "nitrification flux" ;
		F_NIT_vr:units = "gN/m^3/s" ;
		F_NIT_vr:cell_methods = "time: mean" ;
		F_NIT_vr:_FillValue = 1.e+36f ;
		F_NIT_vr:missing_value = 1.e+36f ;
	float GC_HEAT1(time, lndgrid) ;
		GC_HEAT1:long_name = "initial gridcell total heat content" ;
		GC_HEAT1:units = "J/m^2" ;
		GC_HEAT1:cell_methods = "time: mean" ;
		GC_HEAT1:_FillValue = 1.e+36f ;
		GC_HEAT1:missing_value = 1.e+36f ;
	float GC_ICE1(time, lndgrid) ;
		GC_ICE1:long_name = "initial gridcell total ice content" ;
		GC_ICE1:units = "mm" ;
		GC_ICE1:cell_methods = "time: mean" ;
		GC_ICE1:_FillValue = 1.e+36f ;
		GC_ICE1:missing_value = 1.e+36f ;
	float GC_LIQ1(time, lndgrid) ;
		GC_LIQ1:long_name = "initial gridcell total liq content" ;
		GC_LIQ1:units = "mm" ;
		GC_LIQ1:cell_methods = "time: mean" ;
		GC_LIQ1:_FillValue = 1.e+36f ;
		GC_LIQ1:missing_value = 1.e+36f ;
	float GPP(time, lndgrid) ;
		GPP:long_name = "gross primary production" ;
		GPP:units = "gC/m^2/s" ;
		GPP:cell_methods = "time: mean" ;
		GPP:_FillValue = 1.e+36f ;
		GPP:missing_value = 1.e+36f ;
	float GR(time, lndgrid) ;
		GR:long_name = "total growth respiration" ;
		GR:units = "gC/m^2/s" ;
		GR:cell_methods = "time: mean" ;
		GR:_FillValue = 1.e+36f ;
		GR:missing_value = 1.e+36f ;
	float GROSS_NMIN(time, lndgrid) ;
		GROSS_NMIN:long_name = "gross rate of N mineralization" ;
		GROSS_NMIN:units = "gN/m^2/s" ;
		GROSS_NMIN:cell_methods = "time: mean" ;
		GROSS_NMIN:_FillValue = 1.e+36f ;
		GROSS_NMIN:missing_value = 1.e+36f ;
	float H2OCAN(time, lndgrid) ;
		H2OCAN:long_name = "intercepted water" ;
		H2OCAN:units = "mm" ;
		H2OCAN:cell_methods = "time: mean" ;
		H2OCAN:_FillValue = 1.e+36f ;
		H2OCAN:missing_value = 1.e+36f ;
	float H2OSFC(time, lndgrid) ;
		H2OSFC:long_name = "surface water depth" ;
		H2OSFC:units = "mm" ;
		H2OSFC:cell_methods = "time: mean" ;
		H2OSFC:_FillValue = 1.e+36f ;
		H2OSFC:missing_value = 1.e+36f ;
	float H2OSNO(time, lndgrid) ;
		H2OSNO:long_name = "snow depth (liquid water)" ;
		H2OSNO:units = "mm" ;
		H2OSNO:cell_methods = "time: mean" ;
		H2OSNO:_FillValue = 1.e+36f ;
		H2OSNO:missing_value = 1.e+36f ;
	float H2OSNO_TOP(time, lndgrid) ;
		H2OSNO_TOP:long_name = "mass of snow in top snow layer" ;
		H2OSNO_TOP:units = "kg/m2" ;
		H2OSNO_TOP:cell_methods = "time: mean" ;
		H2OSNO_TOP:_FillValue = 1.e+36f ;
		H2OSNO_TOP:missing_value = 1.e+36f ;
	float H2OSOI(time, levgrnd, lndgrid) ;
		H2OSOI:long_name = "volumetric soil water (vegetated landunits only)" ;
		H2OSOI:units = "mm3/mm3" ;
		H2OSOI:cell_methods = "time: mean" ;
		H2OSOI:_FillValue = 1.e+36f ;
		H2OSOI:missing_value = 1.e+36f ;
	float HC(time, lndgrid) ;
		HC:long_name = "heat content of soil/snow/lake" ;
		HC:units = "MJ/m2" ;
		HC:cell_methods = "time: mean" ;
		HC:_FillValue = 1.e+36f ;
		HC:missing_value = 1.e+36f ;
	float HCSOI(time, lndgrid) ;
		HCSOI:long_name = "soil heat content" ;
		HCSOI:units = "MJ/m2" ;
		HCSOI:cell_methods = "time: mean" ;
		HCSOI:_FillValue = 1.e+36f ;
		HCSOI:missing_value = 1.e+36f ;
	float HEAT_FROM_AC(time, lndgrid) ;
		HEAT_FROM_AC:long_name = "sensible heat flux put into canyon due to heat removed from air conditioning" ;
		HEAT_FROM_AC:units = "W/m^2" ;
		HEAT_FROM_AC:cell_methods = "time: mean" ;
		HEAT_FROM_AC:_FillValue = 1.e+36f ;
		HEAT_FROM_AC:missing_value = 1.e+36f ;
	float HR(time, lndgrid) ;
		HR:long_name = "total heterotrophic respiration" ;
		HR:units = "gC/m^2/s" ;
		HR:cell_methods = "time: mean" ;
		HR:_FillValue = 1.e+36f ;
		HR:missing_value = 1.e+36f ;
	float HR_vr(time, levdcmp, lndgrid) ;
		HR_vr:long_name = "total vertically resolved heterotrophic respiration" ;
		HR_vr:units = "gC/m^3/s" ;
		HR_vr:cell_methods = "time: mean" ;
		HR_vr:_FillValue = 1.e+36f ;
		HR_vr:missing_value = 1.e+36f ;
	float HTOP(time, lndgrid) ;
		HTOP:long_name = "canopy top" ;
		HTOP:units = "m" ;
		HTOP:cell_methods = "time: mean" ;
		HTOP:_FillValue = 1.e+36f ;
		HTOP:missing_value = 1.e+36f ;
	float INT_SNOW(time, lndgrid) ;
		INT_SNOW:long_name = "accumulated swe (vegetated landunits only)" ;
		INT_SNOW:units = "mm" ;
		INT_SNOW:cell_methods = "time: mean" ;
		INT_SNOW:_FillValue = 1.e+36f ;
		INT_SNOW:missing_value = 1.e+36f ;
	float LAISHA(time, lndgrid) ;
		LAISHA:long_name = "shaded projected leaf area index" ;
		LAISHA:units = "none" ;
		LAISHA:cell_methods = "time: mean" ;
		LAISHA:_FillValue = 1.e+36f ;
		LAISHA:missing_value = 1.e+36f ;
	float LAISUN(time, lndgrid) ;
		LAISUN:long_name = "sunlit projected leaf area index" ;
		LAISUN:units = "none" ;
		LAISUN:cell_methods = "time: mean" ;
		LAISUN:_FillValue = 1.e+36f ;
		LAISUN:missing_value = 1.e+36f ;
	float LAKEICEFRAC(time, levlak, lndgrid) ;
		LAKEICEFRAC:long_name = "lake layer ice mass fraction" ;
		LAKEICEFRAC:units = "unitless" ;
		LAKEICEFRAC:cell_methods = "time: mean" ;
		LAKEICEFRAC:_FillValue = 1.e+36f ;
		LAKEICEFRAC:missing_value = 1.e+36f ;
	float LAKEICETHICK(time, lndgrid) ;
		LAKEICETHICK:long_name = "thickness of lake ice (including physical expansion on freezing)" ;
		LAKEICETHICK:units = "m" ;
		LAKEICETHICK:cell_methods = "time: mean" ;
		LAKEICETHICK:_FillValue = 1.e+36f ;
		LAKEICETHICK:missing_value = 1.e+36f ;
	float LAND_UPTAKE(time, lndgrid) ;
		LAND_UPTAKE:long_name = "NEE minus LAND_USE_FLUX, negative for update" ;
		LAND_UPTAKE:units = "gC/m^2/s" ;
		LAND_UPTAKE:cell_methods = "time: mean" ;
		LAND_UPTAKE:_FillValue = 1.e+36f ;
		LAND_UPTAKE:missing_value = 1.e+36f ;
	float LAND_USE_FLUX(time, lndgrid) ;
		LAND_USE_FLUX:long_name = "total C emitted from land cover conversion and wood product pools" ;
		LAND_USE_FLUX:units = "gC/m^2/s" ;
		LAND_USE_FLUX:cell_methods = "time: mean" ;
		LAND_USE_FLUX:_FillValue = 1.e+36f ;
		LAND_USE_FLUX:missing_value = 1.e+36f ;
	float LEAFC(time, lndgrid) ;
		LEAFC:long_name = "leaf C" ;
		LEAFC:units = "gC/m^2" ;
		LEAFC:cell_methods = "time: mean" ;
		LEAFC:_FillValue = 1.e+36f ;
		LEAFC:missing_value = 1.e+36f ;
	float LEAFC_ALLOC(time, lndgrid) ;
		LEAFC_ALLOC:long_name = "leaf C allocation" ;
		LEAFC_ALLOC:units = "gC/m^2/s" ;
		LEAFC_ALLOC:cell_methods = "time: mean" ;
		LEAFC_ALLOC:_FillValue = 1.e+36f ;
		LEAFC_ALLOC:missing_value = 1.e+36f ;
	float LEAFC_LOSS(time, lndgrid) ;
		LEAFC_LOSS:long_name = "leaf C loss" ;
		LEAFC_LOSS:units = "gC/m^2/s" ;
		LEAFC_LOSS:cell_methods = "time: mean" ;
		LEAFC_LOSS:_FillValue = 1.e+36f ;
		LEAFC_LOSS:missing_value = 1.e+36f ;
	float LEAFN(time, lndgrid) ;
		LEAFN:long_name = "leaf N" ;
		LEAFN:units = "gN/m^2" ;
		LEAFN:cell_methods = "time: mean" ;
		LEAFN:_FillValue = 1.e+36f ;
		LEAFN:missing_value = 1.e+36f ;
	float LEAF_MR(time, lndgrid) ;
		LEAF_MR:long_name = "leaf maintenance respiration" ;
		LEAF_MR:units = "gC/m^2/s" ;
		LEAF_MR:cell_methods = "time: mean" ;
		LEAF_MR:_FillValue = 1.e+36f ;
		LEAF_MR:missing_value = 1.e+36f ;
	float LFC2(time, lndgrid) ;
		LFC2:long_name = "conversion area fraction of BET and BDT that burned" ;
		LFC2:units = "per sec" ;
		LFC2:cell_methods = "time: mean" ;
		LFC2:_FillValue = 1.e+36f ;
		LFC2:missing_value = 1.e+36f ;
	float LF_CONV_CFLUX(time, lndgrid) ;
		LF_CONV_CFLUX:long_name = "conversion carbon due to BET and BDT area decreasing" ;
		LF_CONV_CFLUX:units = "gC/m^2/s" ;
		LF_CONV_CFLUX:cell_methods = "time: mean" ;
		LF_CONV_CFLUX:_FillValue = 1.e+36f ;
		LF_CONV_CFLUX:missing_value = 1.e+36f ;
	float LITFALL(time, lndgrid) ;
		LITFALL:long_name = "litterfall (leaves and fine roots)" ;
		LITFALL:units = "gC/m^2/s" ;
		LITFALL:cell_methods = "time: mean" ;
		LITFALL:_FillValue = 1.e+36f ;
		LITFALL:missing_value = 1.e+36f ;
	float LITHR(time, lndgrid) ;
		LITHR:long_name = "litter heterotrophic respiration" ;
		LITHR:units = "gC/m^2/s" ;
		LITHR:cell_methods = "time: mean" ;
		LITHR:_FillValue = 1.e+36f ;
		LITHR:missing_value = 1.e+36f ;
	float LITR1C(time, lndgrid) ;
		LITR1C:long_name = "LITR1 C" ;
		LITR1C:units = "gC/m^2" ;
		LITR1C:cell_methods = "time: mean" ;
		LITR1C:_FillValue = 1.e+36f ;
		LITR1C:missing_value = 1.e+36f ;
	float LITR1C_TO_SOIL1C(time, lndgrid) ;
		LITR1C_TO_SOIL1C:long_name = "decomp. of litter 1 C to soil 1 C" ;
		LITR1C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR1C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR1C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR1C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR1C_vr(time, levdcmp, lndgrid) ;
		LITR1C_vr:long_name = "LITR1 C (vertically resolved)" ;
		LITR1C_vr:units = "gC/m^3" ;
		LITR1C_vr:cell_methods = "time: mean" ;
		LITR1C_vr:_FillValue = 1.e+36f ;
		LITR1C_vr:missing_value = 1.e+36f ;
	float LITR1N(time, lndgrid) ;
		LITR1N:long_name = "LITR1 N" ;
		LITR1N:units = "gN/m^2" ;
		LITR1N:cell_methods = "time: mean" ;
		LITR1N:_FillValue = 1.e+36f ;
		LITR1N:missing_value = 1.e+36f ;
	float LITR1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR1N_TNDNCY_VERT_TRANS:long_name = "litter 1 N tendency due to vertical transport" ;
		LITR1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR1N_TO_SOIL1N(time, lndgrid) ;
		LITR1N_TO_SOIL1N:long_name = "decomp. of litter 1 N to soil 1 N" ;
		LITR1N_TO_SOIL1N:units = "gN/m^2" ;
		LITR1N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR1N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR1N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR1N_vr(time, levdcmp, lndgrid) ;
		LITR1N_vr:long_name = "LITR1 N (vertically resolved)" ;
		LITR1N_vr:units = "gN/m^3" ;
		LITR1N_vr:cell_methods = "time: mean" ;
		LITR1N_vr:_FillValue = 1.e+36f ;
		LITR1N_vr:missing_value = 1.e+36f ;
	float LITR1_HR(time, lndgrid) ;
		LITR1_HR:long_name = "Het. Resp. from litter 1" ;
		LITR1_HR:units = "gC/m^2/s" ;
		LITR1_HR:cell_methods = "time: mean" ;
		LITR1_HR:_FillValue = 1.e+36f ;
		LITR1_HR:missing_value = 1.e+36f ;
	float LITR2C(time, lndgrid) ;
		LITR2C:long_name = "LITR2 C" ;
		LITR2C:units = "gC/m^2" ;
		LITR2C:cell_methods = "time: mean" ;
		LITR2C:_FillValue = 1.e+36f ;
		LITR2C:missing_value = 1.e+36f ;
	float LITR2C_TO_SOIL1C(time, lndgrid) ;
		LITR2C_TO_SOIL1C:long_name = "decomp. of litter 2 C to soil 1 C" ;
		LITR2C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR2C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR2C_vr(time, levdcmp, lndgrid) ;
		LITR2C_vr:long_name = "LITR2 C (vertically resolved)" ;
		LITR2C_vr:units = "gC/m^3" ;
		LITR2C_vr:cell_methods = "time: mean" ;
		LITR2C_vr:_FillValue = 1.e+36f ;
		LITR2C_vr:missing_value = 1.e+36f ;
	float LITR2N(time, lndgrid) ;
		LITR2N:long_name = "LITR2 N" ;
		LITR2N:units = "gN/m^2" ;
		LITR2N:cell_methods = "time: mean" ;
		LITR2N:_FillValue = 1.e+36f ;
		LITR2N:missing_value = 1.e+36f ;
	float LITR2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR2N_TNDNCY_VERT_TRANS:long_name = "litter 2 N tendency due to vertical transport" ;
		LITR2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR2N_TO_SOIL1N(time, lndgrid) ;
		LITR2N_TO_SOIL1N:long_name = "decomp. of litter 2 N to soil 1 N" ;
		LITR2N_TO_SOIL1N:units = "gN/m^2" ;
		LITR2N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR2N_vr(time, levdcmp, lndgrid) ;
		LITR2N_vr:long_name = "LITR2 N (vertically resolved)" ;
		LITR2N_vr:units = "gN/m^3" ;
		LITR2N_vr:cell_methods = "time: mean" ;
		LITR2N_vr:_FillValue = 1.e+36f ;
		LITR2N_vr:missing_value = 1.e+36f ;
	float LITR2_HR(time, lndgrid) ;
		LITR2_HR:long_name = "Het. Resp. from litter 2" ;
		LITR2_HR:units = "gC/m^2/s" ;
		LITR2_HR:cell_methods = "time: mean" ;
		LITR2_HR:_FillValue = 1.e+36f ;
		LITR2_HR:missing_value = 1.e+36f ;
	float LITR3C(time, lndgrid) ;
		LITR3C:long_name = "LITR3 C" ;
		LITR3C:units = "gC/m^2" ;
		LITR3C:cell_methods = "time: mean" ;
		LITR3C:_FillValue = 1.e+36f ;
		LITR3C:missing_value = 1.e+36f ;
	float LITR3C_TO_SOIL2C(time, lndgrid) ;
		LITR3C_TO_SOIL2C:long_name = "decomp. of litter 3 C to soil 2 C" ;
		LITR3C_TO_SOIL2C:units = "gC/m^2/s" ;
		LITR3C_TO_SOIL2C:cell_methods = "time: mean" ;
		LITR3C_TO_SOIL2C:_FillValue = 1.e+36f ;
		LITR3C_TO_SOIL2C:missing_value = 1.e+36f ;
	float LITR3C_vr(time, levdcmp, lndgrid) ;
		LITR3C_vr:long_name = "LITR3 C (vertically resolved)" ;
		LITR3C_vr:units = "gC/m^3" ;
		LITR3C_vr:cell_methods = "time: mean" ;
		LITR3C_vr:_FillValue = 1.e+36f ;
		LITR3C_vr:missing_value = 1.e+36f ;
	float LITR3N(time, lndgrid) ;
		LITR3N:long_name = "LITR3 N" ;
		LITR3N:units = "gN/m^2" ;
		LITR3N:cell_methods = "time: mean" ;
		LITR3N:_FillValue = 1.e+36f ;
		LITR3N:missing_value = 1.e+36f ;
	float LITR3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR3N_TNDNCY_VERT_TRANS:long_name = "litter 3 N tendency due to vertical transport" ;
		LITR3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR3N_TO_SOIL2N(time, lndgrid) ;
		LITR3N_TO_SOIL2N:long_name = "decomp. of litter 3 N to soil 2 N" ;
		LITR3N_TO_SOIL2N:units = "gN/m^2" ;
		LITR3N_TO_SOIL2N:cell_methods = "time: mean" ;
		LITR3N_TO_SOIL2N:_FillValue = 1.e+36f ;
		LITR3N_TO_SOIL2N:missing_value = 1.e+36f ;
	float LITR3N_vr(time, levdcmp, lndgrid) ;
		LITR3N_vr:long_name = "LITR3 N (vertically resolved)" ;
		LITR3N_vr:units = "gN/m^3" ;
		LITR3N_vr:cell_methods = "time: mean" ;
		LITR3N_vr:_FillValue = 1.e+36f ;
		LITR3N_vr:missing_value = 1.e+36f ;
	float LITR3_HR(time, lndgrid) ;
		LITR3_HR:long_name = "Het. Resp. from litter 3" ;
		LITR3_HR:units = "gC/m^2/s" ;
		LITR3_HR:cell_methods = "time: mean" ;
		LITR3_HR:_FillValue = 1.e+36f ;
		LITR3_HR:missing_value = 1.e+36f ;
	float LITTERC(time, lndgrid) ;
		LITTERC:long_name = "litter C" ;
		LITTERC:units = "gC/m^2" ;
		LITTERC:cell_methods = "time: mean" ;
		LITTERC:_FillValue = 1.e+36f ;
		LITTERC:missing_value = 1.e+36f ;
	float LITTERC_HR(time, lndgrid) ;
		LITTERC_HR:long_name = "litter C heterotrophic respiration" ;
		LITTERC_HR:units = "gC/m^2/s" ;
		LITTERC_HR:cell_methods = "time: mean" ;
		LITTERC_HR:_FillValue = 1.e+36f ;
		LITTERC_HR:missing_value = 1.e+36f ;
	float LITTERC_LOSS(time, lndgrid) ;
		LITTERC_LOSS:long_name = "litter C loss" ;
		LITTERC_LOSS:units = "gC/m^2/s" ;
		LITTERC_LOSS:cell_methods = "time: mean" ;
		LITTERC_LOSS:_FillValue = 1.e+36f ;
		LITTERC_LOSS:missing_value = 1.e+36f ;
	float LIVECROOTC(time, lndgrid) ;
		LIVECROOTC:long_name = "live coarse root C" ;
		LIVECROOTC:units = "gC/m^2" ;
		LIVECROOTC:cell_methods = "time: mean" ;
		LIVECROOTC:_FillValue = 1.e+36f ;
		LIVECROOTC:missing_value = 1.e+36f ;
	float LIVECROOTN(time, lndgrid) ;
		LIVECROOTN:long_name = "live coarse root N" ;
		LIVECROOTN:units = "gN/m^2" ;
		LIVECROOTN:cell_methods = "time: mean" ;
		LIVECROOTN:_FillValue = 1.e+36f ;
		LIVECROOTN:missing_value = 1.e+36f ;
	float LIVESTEMC(time, lndgrid) ;
		LIVESTEMC:long_name = "live stem C" ;
		LIVESTEMC:units = "gC/m^2" ;
		LIVESTEMC:cell_methods = "time: mean" ;
		LIVESTEMC:_FillValue = 1.e+36f ;
		LIVESTEMC:missing_value = 1.e+36f ;
	float LIVESTEMN(time, lndgrid) ;
		LIVESTEMN:long_name = "live stem N" ;
		LIVESTEMN:units = "gN/m^2" ;
		LIVESTEMN:cell_methods = "time: mean" ;
		LIVESTEMN:_FillValue = 1.e+36f ;
		LIVESTEMN:missing_value = 1.e+36f ;
	float MEG_acetaldehyde(time, lndgrid) ;
		MEG_acetaldehyde:long_name = "MEGAN flux" ;
		MEG_acetaldehyde:units = "kg/m2/sec" ;
		MEG_acetaldehyde:cell_methods = "time: mean" ;
		MEG_acetaldehyde:_FillValue = 1.e+36f ;
		MEG_acetaldehyde:missing_value = 1.e+36f ;
	float MEG_acetic_acid(time, lndgrid) ;
		MEG_acetic_acid:long_name = "MEGAN flux" ;
		MEG_acetic_acid:units = "kg/m2/sec" ;
		MEG_acetic_acid:cell_methods = "time: mean" ;
		MEG_acetic_acid:_FillValue = 1.e+36f ;
		MEG_acetic_acid:missing_value = 1.e+36f ;
	float MEG_acetone(time, lndgrid) ;
		MEG_acetone:long_name = "MEGAN flux" ;
		MEG_acetone:units = "kg/m2/sec" ;
		MEG_acetone:cell_methods = "time: mean" ;
		MEG_acetone:_FillValue = 1.e+36f ;
		MEG_acetone:missing_value = 1.e+36f ;
	float MEG_carene_3(time, lndgrid) ;
		MEG_carene_3:long_name = "MEGAN flux" ;
		MEG_carene_3:units = "kg/m2/sec" ;
		MEG_carene_3:cell_methods = "time: mean" ;
		MEG_carene_3:_FillValue = 1.e+36f ;
		MEG_carene_3:missing_value = 1.e+36f ;
	float MEG_ethanol(time, lndgrid) ;
		MEG_ethanol:long_name = "MEGAN flux" ;
		MEG_ethanol:units = "kg/m2/sec" ;
		MEG_ethanol:cell_methods = "time: mean" ;
		MEG_ethanol:_FillValue = 1.e+36f ;
		MEG_ethanol:missing_value = 1.e+36f ;
	float MEG_formaldehyde(time, lndgrid) ;
		MEG_formaldehyde:long_name = "MEGAN flux" ;
		MEG_formaldehyde:units = "kg/m2/sec" ;
		MEG_formaldehyde:cell_methods = "time: mean" ;
		MEG_formaldehyde:_FillValue = 1.e+36f ;
		MEG_formaldehyde:missing_value = 1.e+36f ;
	float MEG_isoprene(time, lndgrid) ;
		MEG_isoprene:long_name = "MEGAN flux" ;
		MEG_isoprene:units = "kg/m2/sec" ;
		MEG_isoprene:cell_methods = "time: mean" ;
		MEG_isoprene:_FillValue = 1.e+36f ;
		MEG_isoprene:missing_value = 1.e+36f ;
	float MEG_methanol(time, lndgrid) ;
		MEG_methanol:long_name = "MEGAN flux" ;
		MEG_methanol:units = "kg/m2/sec" ;
		MEG_methanol:cell_methods = "time: mean" ;
		MEG_methanol:_FillValue = 1.e+36f ;
		MEG_methanol:missing_value = 1.e+36f ;
	float MEG_pinene_a(time, lndgrid) ;
		MEG_pinene_a:long_name = "MEGAN flux" ;
		MEG_pinene_a:units = "kg/m2/sec" ;
		MEG_pinene_a:cell_methods = "time: mean" ;
		MEG_pinene_a:_FillValue = 1.e+36f ;
		MEG_pinene_a:missing_value = 1.e+36f ;
	float MEG_thujene_a(time, lndgrid) ;
		MEG_thujene_a:long_name = "MEGAN flux" ;
		MEG_thujene_a:units = "kg/m2/sec" ;
		MEG_thujene_a:cell_methods = "time: mean" ;
		MEG_thujene_a:_FillValue = 1.e+36f ;
		MEG_thujene_a:missing_value = 1.e+36f ;
	float MR(time, lndgrid) ;
		MR:long_name = "maintenance respiration" ;
		MR:units = "gC/m^2/s" ;
		MR:cell_methods = "time: mean" ;
		MR:_FillValue = 1.e+36f ;
		MR:missing_value = 1.e+36f ;
	float M_LITR1C_TO_LEACHING(time, lndgrid) ;
		M_LITR1C_TO_LEACHING:long_name = "litter 1 C leaching loss" ;
		M_LITR1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR2C_TO_LEACHING(time, lndgrid) ;
		M_LITR2C_TO_LEACHING:long_name = "litter 2 C leaching loss" ;
		M_LITR2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR3C_TO_LEACHING(time, lndgrid) ;
		M_LITR3C_TO_LEACHING:long_name = "litter 3 C leaching loss" ;
		M_LITR3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR3C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL1C_TO_LEACHING(time, lndgrid) ;
		M_SOIL1C_TO_LEACHING:long_name = "soil 1 C leaching loss" ;
		M_SOIL1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL2C_TO_LEACHING(time, lndgrid) ;
		M_SOIL2C_TO_LEACHING:long_name = "soil 2 C leaching loss" ;
		M_SOIL2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL3C_TO_LEACHING(time, lndgrid) ;
		M_SOIL3C_TO_LEACHING:long_name = "soil 3 C leaching loss" ;
		M_SOIL3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL3C_TO_LEACHING:missing_value = 1.e+36f ;
	float NBP(time, lndgrid) ;
		NBP:long_name = "net biome production, includes fire, landuse, and harvest flux, positive for sink" ;
		NBP:units = "gC/m^2/s" ;
		NBP:cell_methods = "time: mean" ;
		NBP:_FillValue = 1.e+36f ;
		NBP:missing_value = 1.e+36f ;
	float NDEPLOY(time, lndgrid) ;
		NDEPLOY:long_name = "total N deployed in new growth" ;
		NDEPLOY:units = "gN/m^2/s" ;
		NDEPLOY:cell_methods = "time: mean" ;
		NDEPLOY:_FillValue = 1.e+36f ;
		NDEPLOY:missing_value = 1.e+36f ;
	float NDEP_TO_SMINN(time, lndgrid) ;
		NDEP_TO_SMINN:long_name = "atmospheric N deposition to soil mineral N" ;
		NDEP_TO_SMINN:units = "gN/m^2/s" ;
		NDEP_TO_SMINN:cell_methods = "time: mean" ;
		NDEP_TO_SMINN:_FillValue = 1.e+36f ;
		NDEP_TO_SMINN:missing_value = 1.e+36f ;
	float NEE(time, lndgrid) ;
		NEE:long_name = "net ecosystem exchange of carbon, includes fire, landuse, harvest, and hrv_xsmrpool flux, positive for source" ;
		NEE:units = "gC/m^2/s" ;
		NEE:cell_methods = "time: mean" ;
		NEE:_FillValue = 1.e+36f ;
		NEE:missing_value = 1.e+36f ;
	float NEM(time, lndgrid) ;
		NEM:long_name = "Gridcell net adjustment to NEE passed to atm. for methane production" ;
		NEM:units = "gC/m2/s" ;
		NEM:cell_methods = "time: mean" ;
		NEM:_FillValue = 1.e+36f ;
		NEM:missing_value = 1.e+36f ;
	float NEP(time, lndgrid) ;
		NEP:long_name = "net ecosystem production, excludes fire, landuse, and harvest flux, positive for sink" ;
		NEP:units = "gC/m^2/s" ;
		NEP:cell_methods = "time: mean" ;
		NEP:_FillValue = 1.e+36f ;
		NEP:missing_value = 1.e+36f ;
	float NET_NMIN(time, lndgrid) ;
		NET_NMIN:long_name = "net rate of N mineralization" ;
		NET_NMIN:units = "gN/m^2/s" ;
		NET_NMIN:cell_methods = "time: mean" ;
		NET_NMIN:_FillValue = 1.e+36f ;
		NET_NMIN:missing_value = 1.e+36f ;
	float NFIRE(time, lndgrid) ;
		NFIRE:long_name = "fire counts valid only in Reg.C" ;
		NFIRE:units = "counts/km2/sec" ;
		NFIRE:cell_methods = "time: mean" ;
		NFIRE:_FillValue = 1.e+36f ;
		NFIRE:missing_value = 1.e+36f ;
	float NFIX_TO_SMINN(time, lndgrid) ;
		NFIX_TO_SMINN:long_name = "symbiotic/asymbiotic N fixation to soil mineral N" ;
		NFIX_TO_SMINN:units = "gN/m^2/s" ;
		NFIX_TO_SMINN:cell_methods = "time: mean" ;
		NFIX_TO_SMINN:_FillValue = 1.e+36f ;
		NFIX_TO_SMINN:missing_value = 1.e+36f ;
	float NPP(time, lndgrid) ;
		NPP:long_name = "net primary production" ;
		NPP:units = "gC/m^2/s" ;
		NPP:cell_methods = "time: mean" ;
		NPP:_FillValue = 1.e+36f ;
		NPP:missing_value = 1.e+36f ;
	float OCDEP(time, lndgrid) ;
		OCDEP:long_name = "total OC deposition (dry+wet) from atmosphere" ;
		OCDEP:units = "kg/m^2/s" ;
		OCDEP:cell_methods = "time: mean" ;
		OCDEP:_FillValue = 1.e+36f ;
		OCDEP:missing_value = 1.e+36f ;
	float O_SCALAR(time, levdcmp, lndgrid) ;
		O_SCALAR:long_name = "fraction by which decomposition is reduced due to anoxia" ;
		O_SCALAR:units = "unitless" ;
		O_SCALAR:cell_methods = "time: mean" ;
		O_SCALAR:_FillValue = 1.e+36f ;
		O_SCALAR:missing_value = 1.e+36f ;
	float PARVEGLN(time, lndgrid) ;
		PARVEGLN:long_name = "absorbed par by vegetation at local noon" ;
		PARVEGLN:units = "W/m^2" ;
		PARVEGLN:cell_methods = "time: mean" ;
		PARVEGLN:_FillValue = 1.e+36f ;
		PARVEGLN:missing_value = 1.e+36f ;
	float PBOT(time, lndgrid) ;
		PBOT:long_name = "atmospheric pressure" ;
		PBOT:units = "Pa" ;
		PBOT:cell_methods = "time: mean" ;
		PBOT:_FillValue = 1.e+36f ;
		PBOT:missing_value = 1.e+36f ;
	float PCH4(time, lndgrid) ;
		PCH4:long_name = "atmospheric partial pressure of CH4" ;
		PCH4:units = "Pa" ;
		PCH4:cell_methods = "time: mean" ;
		PCH4:_FillValue = 1.e+36f ;
		PCH4:missing_value = 1.e+36f ;
	float PCO2(time, lndgrid) ;
		PCO2:long_name = "atmospheric partial pressure of CO2" ;
		PCO2:units = "Pa" ;
		PCO2:cell_methods = "time: mean" ;
		PCO2:_FillValue = 1.e+36f ;
		PCO2:missing_value = 1.e+36f ;
	float PCT_LANDUNIT(time, ltype, lndgrid) ;
		PCT_LANDUNIT:long_name = "% of each landunit on grid cell" ;
		PCT_LANDUNIT:units = "%" ;
		PCT_LANDUNIT:cell_methods = "time: mean" ;
		PCT_LANDUNIT:_FillValue = 1.e+36f ;
		PCT_LANDUNIT:missing_value = 1.e+36f ;
	float PCT_NAT_PFT(time, natpft, lndgrid) ;
		PCT_NAT_PFT:long_name = "% of each PFT on the natural vegetation (i.e., soil) landunit" ;
		PCT_NAT_PFT:units = "%" ;
		PCT_NAT_PFT:cell_methods = "time: mean" ;
		PCT_NAT_PFT:_FillValue = 1.e+36f ;
		PCT_NAT_PFT:missing_value = 1.e+36f ;
	float PFT_CTRUNC(time, lndgrid) ;
		PFT_CTRUNC:long_name = "pft-level sink for C truncation" ;
		PFT_CTRUNC:units = "gC/m^2" ;
		PFT_CTRUNC:cell_methods = "time: mean" ;
		PFT_CTRUNC:_FillValue = 1.e+36f ;
		PFT_CTRUNC:missing_value = 1.e+36f ;
	float PFT_FIRE_CLOSS(time, lndgrid) ;
		PFT_FIRE_CLOSS:long_name = "total pft-level fire C loss for non-peat fires outside land-type converted region" ;
		PFT_FIRE_CLOSS:units = "gC/m^2/s" ;
		PFT_FIRE_CLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_CLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_CLOSS:missing_value = 1.e+36f ;
	float PFT_FIRE_NLOSS(time, lndgrid) ;
		PFT_FIRE_NLOSS:long_name = "total pft-level fire N loss" ;
		PFT_FIRE_NLOSS:units = "gN/m^2/s" ;
		PFT_FIRE_NLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_NLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_NLOSS:missing_value = 1.e+36f ;
	float PFT_NTRUNC(time, lndgrid) ;
		PFT_NTRUNC:long_name = "pft-level sink for N truncation" ;
		PFT_NTRUNC:units = "gN/m^2" ;
		PFT_NTRUNC:cell_methods = "time: mean" ;
		PFT_NTRUNC:_FillValue = 1.e+36f ;
		PFT_NTRUNC:missing_value = 1.e+36f ;
	float PLANT_NDEMAND(time, lndgrid) ;
		PLANT_NDEMAND:long_name = "N flux required to support initial GPP" ;
		PLANT_NDEMAND:units = "gN/m^2/s" ;
		PLANT_NDEMAND:cell_methods = "time: mean" ;
		PLANT_NDEMAND:_FillValue = 1.e+36f ;
		PLANT_NDEMAND:missing_value = 1.e+36f ;
	float POTENTIAL_IMMOB(time, lndgrid) ;
		POTENTIAL_IMMOB:long_name = "potential N immobilization" ;
		POTENTIAL_IMMOB:units = "gN/m^2/s" ;
		POTENTIAL_IMMOB:cell_methods = "time: mean" ;
		POTENTIAL_IMMOB:_FillValue = 1.e+36f ;
		POTENTIAL_IMMOB:missing_value = 1.e+36f ;
	float POT_F_DENIT(time, lndgrid) ;
		POT_F_DENIT:long_name = "potential denitrification flux" ;
		POT_F_DENIT:units = "gN/m^2/s" ;
		POT_F_DENIT:cell_methods = "time: mean" ;
		POT_F_DENIT:_FillValue = 1.e+36f ;
		POT_F_DENIT:missing_value = 1.e+36f ;
	float POT_F_NIT(time, lndgrid) ;
		POT_F_NIT:long_name = "potential nitrification flux" ;
		POT_F_NIT:units = "gN/m^2/s" ;
		POT_F_NIT:cell_methods = "time: mean" ;
		POT_F_NIT:_FillValue = 1.e+36f ;
		POT_F_NIT:missing_value = 1.e+36f ;
	float PROD100C(time, lndgrid) ;
		PROD100C:long_name = "100-yr wood product C" ;
		PROD100C:units = "gC/m^2" ;
		PROD100C:cell_methods = "time: mean" ;
		PROD100C:_FillValue = 1.e+36f ;
		PROD100C:missing_value = 1.e+36f ;
	float PROD100C_LOSS(time, lndgrid) ;
		PROD100C_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100C_LOSS:units = "gC/m^2/s" ;
		PROD100C_LOSS:cell_methods = "time: mean" ;
		PROD100C_LOSS:_FillValue = 1.e+36f ;
		PROD100C_LOSS:missing_value = 1.e+36f ;
	float PROD100N(time, lndgrid) ;
		PROD100N:long_name = "100-yr wood product N" ;
		PROD100N:units = "gN/m^2" ;
		PROD100N:cell_methods = "time: mean" ;
		PROD100N:_FillValue = 1.e+36f ;
		PROD100N:missing_value = 1.e+36f ;
	float PROD100N_LOSS(time, lndgrid) ;
		PROD100N_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100N_LOSS:units = "gN/m^2/s" ;
		PROD100N_LOSS:cell_methods = "time: mean" ;
		PROD100N_LOSS:_FillValue = 1.e+36f ;
		PROD100N_LOSS:missing_value = 1.e+36f ;
	float PROD10C(time, lndgrid) ;
		PROD10C:long_name = "10-yr wood product C" ;
		PROD10C:units = "gC/m^2" ;
		PROD10C:cell_methods = "time: mean" ;
		PROD10C:_FillValue = 1.e+36f ;
		PROD10C:missing_value = 1.e+36f ;
	float PROD10C_LOSS(time, lndgrid) ;
		PROD10C_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10C_LOSS:units = "gC/m^2/s" ;
		PROD10C_LOSS:cell_methods = "time: mean" ;
		PROD10C_LOSS:_FillValue = 1.e+36f ;
		PROD10C_LOSS:missing_value = 1.e+36f ;
	float PROD10N(time, lndgrid) ;
		PROD10N:long_name = "10-yr wood product N" ;
		PROD10N:units = "gN/m^2" ;
		PROD10N:cell_methods = "time: mean" ;
		PROD10N:_FillValue = 1.e+36f ;
		PROD10N:missing_value = 1.e+36f ;
	float PROD10N_LOSS(time, lndgrid) ;
		PROD10N_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10N_LOSS:units = "gN/m^2/s" ;
		PROD10N_LOSS:cell_methods = "time: mean" ;
		PROD10N_LOSS:_FillValue = 1.e+36f ;
		PROD10N_LOSS:missing_value = 1.e+36f ;
	float PRODUCT_CLOSS(time, lndgrid) ;
		PRODUCT_CLOSS:long_name = "total carbon loss from wood product pools" ;
		PRODUCT_CLOSS:units = "gC/m^2/s" ;
		PRODUCT_CLOSS:cell_methods = "time: mean" ;
		PRODUCT_CLOSS:_FillValue = 1.e+36f ;
		PRODUCT_CLOSS:missing_value = 1.e+36f ;
	float PRODUCT_NLOSS(time, lndgrid) ;
		PRODUCT_NLOSS:long_name = "total N loss from wood product pools" ;
		PRODUCT_NLOSS:units = "gN/m^2/s" ;
		PRODUCT_NLOSS:cell_methods = "time: mean" ;
		PRODUCT_NLOSS:_FillValue = 1.e+36f ;
		PRODUCT_NLOSS:missing_value = 1.e+36f ;
	float PSNSHA(time, lndgrid) ;
		PSNSHA:long_name = "shaded leaf photosynthesis" ;
		PSNSHA:units = "umolCO2/m^2/s" ;
		PSNSHA:cell_methods = "time: mean" ;
		PSNSHA:_FillValue = 1.e+36f ;
		PSNSHA:missing_value = 1.e+36f ;
	float PSNSHADE_TO_CPOOL(time, lndgrid) ;
		PSNSHADE_TO_CPOOL:long_name = "C fixation from shaded canopy" ;
		PSNSHADE_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSHADE_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSHADE_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSHADE_TO_CPOOL:missing_value = 1.e+36f ;
	float PSNSUN(time, lndgrid) ;
		PSNSUN:long_name = "sunlit leaf photosynthesis" ;
		PSNSUN:units = "umolCO2/m^2/s" ;
		PSNSUN:cell_methods = "time: mean" ;
		PSNSUN:_FillValue = 1.e+36f ;
		PSNSUN:missing_value = 1.e+36f ;
	float PSNSUN_TO_CPOOL(time, lndgrid) ;
		PSNSUN_TO_CPOOL:long_name = "C fixation from sunlit canopy" ;
		PSNSUN_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSUN_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSUN_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSUN_TO_CPOOL:missing_value = 1.e+36f ;
	float Q2M(time, lndgrid) ;
		Q2M:long_name = "2m specific humidity" ;
		Q2M:units = "kg/kg" ;
		Q2M:cell_methods = "time: mean" ;
		Q2M:_FillValue = 1.e+36f ;
		Q2M:missing_value = 1.e+36f ;
	float QBOT(time, lndgrid) ;
		QBOT:long_name = "atmospheric specific humidity" ;
		QBOT:units = "kg/kg" ;
		QBOT:cell_methods = "time: mean" ;
		QBOT:_FillValue = 1.e+36f ;
		QBOT:missing_value = 1.e+36f ;
	float QCHARGE(time, lndgrid) ;
		QCHARGE:long_name = "aquifer recharge rate (vegetated landunits only)" ;
		QCHARGE:units = "mm/s" ;
		QCHARGE:cell_methods = "time: mean" ;
		QCHARGE:_FillValue = 1.e+36f ;
		QCHARGE:missing_value = 1.e+36f ;
	float QDRAI(time, lndgrid) ;
		QDRAI:long_name = "sub-surface drainage" ;
		QDRAI:units = "mm/s" ;
		QDRAI:cell_methods = "time: mean" ;
		QDRAI:_FillValue = 1.e+36f ;
		QDRAI:missing_value = 1.e+36f ;
	float QDRAI_PERCH(time, lndgrid) ;
		QDRAI_PERCH:long_name = "perched wt drainage" ;
		QDRAI_PERCH:units = "mm/s" ;
		QDRAI_PERCH:cell_methods = "time: mean" ;
		QDRAI_PERCH:_FillValue = 1.e+36f ;
		QDRAI_PERCH:missing_value = 1.e+36f ;
	float QDRAI_XS(time, lndgrid) ;
		QDRAI_XS:long_name = "saturation excess drainage" ;
		QDRAI_XS:units = "mm/s" ;
		QDRAI_XS:cell_methods = "time: mean" ;
		QDRAI_XS:_FillValue = 1.e+36f ;
		QDRAI_XS:missing_value = 1.e+36f ;
	float QDRIP(time, lndgrid) ;
		QDRIP:long_name = "throughfall" ;
		QDRIP:units = "mm/s" ;
		QDRIP:cell_methods = "time: mean" ;
		QDRIP:_FillValue = 1.e+36f ;
		QDRIP:missing_value = 1.e+36f ;
	float QFLOOD(time, lndgrid) ;
		QFLOOD:long_name = "runoff from river flooding" ;
		QFLOOD:units = "mm/s" ;
		QFLOOD:cell_methods = "time: mean" ;
		QFLOOD:_FillValue = 1.e+36f ;
		QFLOOD:missing_value = 1.e+36f ;
	float QFLX_ICE_DYNBAL(time, lndgrid) ;
		QFLX_ICE_DYNBAL:long_name = "ice dynamic land cover change conversion runoff flux" ;
		QFLX_ICE_DYNBAL:units = "mm/s" ;
		QFLX_ICE_DYNBAL:cell_methods = "time: mean" ;
		QFLX_ICE_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_ICE_DYNBAL:missing_value = 1.e+36f ;
	float QFLX_LIQ_DYNBAL(time, lndgrid) ;
		QFLX_LIQ_DYNBAL:long_name = "liq dynamic land cover change conversion runoff flux" ;
		QFLX_LIQ_DYNBAL:units = "mm/s" ;
		QFLX_LIQ_DYNBAL:cell_methods = "time: mean" ;
		QFLX_LIQ_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_LIQ_DYNBAL:missing_value = 1.e+36f ;
	float QH2OSFC(time, lndgrid) ;
		QH2OSFC:long_name = "surface water runoff" ;
		QH2OSFC:units = "mm/s" ;
		QH2OSFC:cell_methods = "time: mean" ;
		QH2OSFC:_FillValue = 1.e+36f ;
		QH2OSFC:missing_value = 1.e+36f ;
	float QINFL(time, lndgrid) ;
		QINFL:long_name = "infiltration" ;
		QINFL:units = "mm/s" ;
		QINFL:cell_methods = "time: mean" ;
		QINFL:_FillValue = 1.e+36f ;
		QINFL:missing_value = 1.e+36f ;
	float QINTR(time, lndgrid) ;
		QINTR:long_name = "interception" ;
		QINTR:units = "mm/s" ;
		QINTR:cell_methods = "time: mean" ;
		QINTR:_FillValue = 1.e+36f ;
		QINTR:missing_value = 1.e+36f ;
	float QIRRIG(time, lndgrid) ;
		QIRRIG:long_name = "water added through irrigation" ;
		QIRRIG:units = "mm/s" ;
		QIRRIG:cell_methods = "time: mean" ;
		QIRRIG:_FillValue = 1.e+36f ;
		QIRRIG:missing_value = 1.e+36f ;
	float QOVER(time, lndgrid) ;
		QOVER:long_name = "surface runoff" ;
		QOVER:units = "mm/s" ;
		QOVER:cell_methods = "time: mean" ;
		QOVER:_FillValue = 1.e+36f ;
		QOVER:missing_value = 1.e+36f ;
	float QOVER_LAG(time, lndgrid) ;
		QOVER_LAG:long_name = "time-lagged surface runoff for soil columns" ;
		QOVER_LAG:units = "mm/s" ;
		QOVER_LAG:cell_methods = "time: mean" ;
		QOVER_LAG:_FillValue = 1.e+36f ;
		QOVER_LAG:missing_value = 1.e+36f ;
	float QRGWL(time, lndgrid) ;
		QRGWL:long_name = "surface runoff at glaciers (liquid only), wetlands, lakes" ;
		QRGWL:units = "mm/s" ;
		QRGWL:cell_methods = "time: mean" ;
		QRGWL:_FillValue = 1.e+36f ;
		QRGWL:missing_value = 1.e+36f ;
	float QRUNOFF(time, lndgrid) ;
		QRUNOFF:long_name = "total liquid runoff (does not include QSNWCPICE)" ;
		QRUNOFF:units = "mm/s" ;
		QRUNOFF:cell_methods = "time: mean" ;
		QRUNOFF:_FillValue = 1.e+36f ;
		QRUNOFF:missing_value = 1.e+36f ;
	float QRUNOFF_NODYNLNDUSE(time, lndgrid) ;
		QRUNOFF_NODYNLNDUSE:long_name = "total liquid runoff (does not include QSNWCPICE) not including correction for land use change" ;
		QRUNOFF_NODYNLNDUSE:units = "mm/s" ;
		QRUNOFF_NODYNLNDUSE:cell_methods = "time: mean" ;
		QRUNOFF_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QRUNOFF_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QRUNOFF_R(time, lndgrid) ;
		QRUNOFF_R:long_name = "Rural total runoff" ;
		QRUNOFF_R:units = "mm/s" ;
		QRUNOFF_R:cell_methods = "time: mean" ;
		QRUNOFF_R:_FillValue = 1.e+36f ;
		QRUNOFF_R:missing_value = 1.e+36f ;
	float QRUNOFF_U(time, lndgrid) ;
		QRUNOFF_U:long_name = "Urban total runoff" ;
		QRUNOFF_U:units = "mm/s" ;
		QRUNOFF_U:cell_methods = "time: mean" ;
		QRUNOFF_U:_FillValue = 1.e+36f ;
		QRUNOFF_U:missing_value = 1.e+36f ;
	float QSNOMELT(time, lndgrid) ;
		QSNOMELT:long_name = "snow melt" ;
		QSNOMELT:units = "mm/s" ;
		QSNOMELT:cell_methods = "time: mean" ;
		QSNOMELT:_FillValue = 1.e+36f ;
		QSNOMELT:missing_value = 1.e+36f ;
	float QSNWCPICE(time, lndgrid) ;
		QSNWCPICE:long_name = "excess snowfall due to snow capping" ;
		QSNWCPICE:units = "mm/s" ;
		QSNWCPICE:cell_methods = "time: mean" ;
		QSNWCPICE:_FillValue = 1.e+36f ;
		QSNWCPICE:missing_value = 1.e+36f ;
	float QSNWCPICE_NODYNLNDUSE(time, lndgrid) ;
		QSNWCPICE_NODYNLNDUSE:long_name = "excess snowfall due to snow capping not including correction for land use change" ;
		QSNWCPICE_NODYNLNDUSE:units = "mm H2O/s" ;
		QSNWCPICE_NODYNLNDUSE:cell_methods = "time: mean" ;
		QSNWCPICE_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QSNWCPICE_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QSOIL(time, lndgrid) ;
		QSOIL:long_name = "Ground evaporation (soil/snow evaporation + soil/snow sublimation - dew)" ;
		QSOIL:units = "mm/s" ;
		QSOIL:cell_methods = "time: mean" ;
		QSOIL:_FillValue = 1.e+36f ;
		QSOIL:missing_value = 1.e+36f ;
	float QVEGE(time, lndgrid) ;
		QVEGE:long_name = "canopy evaporation" ;
		QVEGE:units = "mm/s" ;
		QVEGE:cell_methods = "time: mean" ;
		QVEGE:_FillValue = 1.e+36f ;
		QVEGE:missing_value = 1.e+36f ;
	float QVEGT(time, lndgrid) ;
		QVEGT:long_name = "canopy transpiration" ;
		QVEGT:units = "mm/s" ;
		QVEGT:cell_methods = "time: mean" ;
		QVEGT:_FillValue = 1.e+36f ;
		QVEGT:missing_value = 1.e+36f ;
	float RAIN(time, lndgrid) ;
		RAIN:long_name = "atmospheric rain" ;
		RAIN:units = "mm/s" ;
		RAIN:cell_methods = "time: mean" ;
		RAIN:_FillValue = 1.e+36f ;
		RAIN:missing_value = 1.e+36f ;
	float RETRANSN(time, lndgrid) ;
		RETRANSN:long_name = "plant pool of retranslocated N" ;
		RETRANSN:units = "gN/m^2" ;
		RETRANSN:cell_methods = "time: mean" ;
		RETRANSN:_FillValue = 1.e+36f ;
		RETRANSN:missing_value = 1.e+36f ;
	float RETRANSN_TO_NPOOL(time, lndgrid) ;
		RETRANSN_TO_NPOOL:long_name = "deployment of retranslocated N" ;
		RETRANSN_TO_NPOOL:units = "gN/m^2/s" ;
		RETRANSN_TO_NPOOL:cell_methods = "time: mean" ;
		RETRANSN_TO_NPOOL:_FillValue = 1.e+36f ;
		RETRANSN_TO_NPOOL:missing_value = 1.e+36f ;
	float RH2M(time, lndgrid) ;
		RH2M:long_name = "2m relative humidity" ;
		RH2M:units = "%" ;
		RH2M:cell_methods = "time: mean" ;
		RH2M:_FillValue = 1.e+36f ;
		RH2M:missing_value = 1.e+36f ;
	float RH2M_R(time, lndgrid) ;
		RH2M_R:long_name = "Rural 2m specific humidity" ;
		RH2M_R:units = "%" ;
		RH2M_R:cell_methods = "time: mean" ;
		RH2M_R:_FillValue = 1.e+36f ;
		RH2M_R:missing_value = 1.e+36f ;
	float RH2M_U(time, lndgrid) ;
		RH2M_U:long_name = "Urban 2m relative humidity" ;
		RH2M_U:units = "%" ;
		RH2M_U:cell_methods = "time: mean" ;
		RH2M_U:_FillValue = 1.e+36f ;
		RH2M_U:missing_value = 1.e+36f ;
	float RR(time, lndgrid) ;
		RR:long_name = "root respiration (fine root MR + total root GR)" ;
		RR:units = "gC/m^2/s" ;
		RR:cell_methods = "time: mean" ;
		RR:_FillValue = 1.e+36f ;
		RR:missing_value = 1.e+36f ;
	float SABG(time, lndgrid) ;
		SABG:long_name = "solar rad absorbed by ground" ;
		SABG:units = "W/m^2" ;
		SABG:cell_methods = "time: mean" ;
		SABG:_FillValue = 1.e+36f ;
		SABG:missing_value = 1.e+36f ;
	float SABG_PEN(time, lndgrid) ;
		SABG_PEN:long_name = "Rural solar rad penetrating top soil or snow layer" ;
		SABG_PEN:units = "watt/m^2" ;
		SABG_PEN:cell_methods = "time: mean" ;
		SABG_PEN:_FillValue = 1.e+36f ;
		SABG_PEN:missing_value = 1.e+36f ;
	float SABV(time, lndgrid) ;
		SABV:long_name = "solar rad absorbed by veg" ;
		SABV:units = "W/m^2" ;
		SABV:cell_methods = "time: mean" ;
		SABV:_FillValue = 1.e+36f ;
		SABV:missing_value = 1.e+36f ;
	float SEEDC(time, lndgrid) ;
		SEEDC:long_name = "pool for seeding new PFTs" ;
		SEEDC:units = "gC/m^2" ;
		SEEDC:cell_methods = "time: mean" ;
		SEEDC:_FillValue = 1.e+36f ;
		SEEDC:missing_value = 1.e+36f ;
	float SEEDN(time, lndgrid) ;
		SEEDN:long_name = "pool for seeding new PFTs" ;
		SEEDN:units = "gN/m^2" ;
		SEEDN:cell_methods = "time: mean" ;
		SEEDN:_FillValue = 1.e+36f ;
		SEEDN:missing_value = 1.e+36f ;
	float SMINN(time, lndgrid) ;
		SMINN:long_name = "soil mineral N" ;
		SMINN:units = "gN/m^2" ;
		SMINN:cell_methods = "time: mean" ;
		SMINN:_FillValue = 1.e+36f ;
		SMINN:missing_value = 1.e+36f ;
	float SMINN_TO_NPOOL(time, lndgrid) ;
		SMINN_TO_NPOOL:long_name = "deployment of soil mineral N uptake" ;
		SMINN_TO_NPOOL:units = "gN/m^2/s" ;
		SMINN_TO_NPOOL:cell_methods = "time: mean" ;
		SMINN_TO_NPOOL:_FillValue = 1.e+36f ;
		SMINN_TO_NPOOL:missing_value = 1.e+36f ;
	float SMINN_TO_PLANT(time, lndgrid) ;
		SMINN_TO_PLANT:long_name = "plant uptake of soil mineral N" ;
		SMINN_TO_PLANT:units = "gN/m^2/s" ;
		SMINN_TO_PLANT:cell_methods = "time: mean" ;
		SMINN_TO_PLANT:_FillValue = 1.e+36f ;
		SMINN_TO_PLANT:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L1(time, lndgrid) ;
		SMINN_TO_SOIL1N_L1:long_name = "mineral N flux for decomp. of LITR1to SOIL1" ;
		SMINN_TO_SOIL1N_L1:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L2(time, lndgrid) ;
		SMINN_TO_SOIL1N_L2:long_name = "mineral N flux for decomp. of LITR2to SOIL1" ;
		SMINN_TO_SOIL1N_L2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S2(time, lndgrid) ;
		SMINN_TO_SOIL1N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL1" ;
		SMINN_TO_SOIL1N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S3(time, lndgrid) ;
		SMINN_TO_SOIL1N_S3:long_name = "mineral N flux for decomp. of SOIL3to SOIL1" ;
		SMINN_TO_SOIL1N_S3:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_L3(time, lndgrid) ;
		SMINN_TO_SOIL2N_L3:long_name = "mineral N flux for decomp. of LITR3to SOIL2" ;
		SMINN_TO_SOIL2N_L3:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_L3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_L3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_L3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_S1(time, lndgrid) ;
		SMINN_TO_SOIL2N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL2" ;
		SMINN_TO_SOIL2N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S1(time, lndgrid) ;
		SMINN_TO_SOIL3N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL3" ;
		SMINN_TO_SOIL3N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S2(time, lndgrid) ;
		SMINN_TO_SOIL3N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL3" ;
		SMINN_TO_SOIL3N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S2:missing_value = 1.e+36f ;
	float SMIN_NH4(time, lndgrid) ;
		SMIN_NH4:long_name = "soil mineral NH4" ;
		SMIN_NH4:units = "gN/m^2" ;
		SMIN_NH4:cell_methods = "time: mean" ;
		SMIN_NH4:_FillValue = 1.e+36f ;
		SMIN_NH4:missing_value = 1.e+36f ;
	float SMIN_NH4_vr(time, levdcmp, lndgrid) ;
		SMIN_NH4_vr:long_name = "soil mineral NH4 (vert. res.)" ;
		SMIN_NH4_vr:units = "gN/m^3" ;
		SMIN_NH4_vr:cell_methods = "time: mean" ;
		SMIN_NH4_vr:_FillValue = 1.e+36f ;
		SMIN_NH4_vr:missing_value = 1.e+36f ;
	float SMIN_NO3(time, lndgrid) ;
		SMIN_NO3:long_name = "soil mineral NO3" ;
		SMIN_NO3:units = "gN/m^2" ;
		SMIN_NO3:cell_methods = "time: mean" ;
		SMIN_NO3:_FillValue = 1.e+36f ;
		SMIN_NO3:missing_value = 1.e+36f ;
	float SMIN_NO3_LEACHED(time, lndgrid) ;
		SMIN_NO3_LEACHED:long_name = "soil NO3 pool loss to leaching" ;
		SMIN_NO3_LEACHED:units = "gN/m^2/s" ;
		SMIN_NO3_LEACHED:cell_methods = "time: mean" ;
		SMIN_NO3_LEACHED:_FillValue = 1.e+36f ;
		SMIN_NO3_LEACHED:missing_value = 1.e+36f ;
	float SMIN_NO3_RUNOFF(time, lndgrid) ;
		SMIN_NO3_RUNOFF:long_name = "soil NO3 pool loss to runoff" ;
		SMIN_NO3_RUNOFF:units = "gN/m^2/s" ;
		SMIN_NO3_RUNOFF:cell_methods = "time: mean" ;
		SMIN_NO3_RUNOFF:_FillValue = 1.e+36f ;
		SMIN_NO3_RUNOFF:missing_value = 1.e+36f ;
	float SMIN_NO3_vr(time, levdcmp, lndgrid) ;
		SMIN_NO3_vr:long_name = "soil mineral NO3 (vert. res.)" ;
		SMIN_NO3_vr:units = "gN/m^3" ;
		SMIN_NO3_vr:cell_methods = "time: mean" ;
		SMIN_NO3_vr:_FillValue = 1.e+36f ;
		SMIN_NO3_vr:missing_value = 1.e+36f ;
	float SNOBCMCL(time, lndgrid) ;
		SNOBCMCL:long_name = "mass of BC in snow column" ;
		SNOBCMCL:units = "kg/m2" ;
		SNOBCMCL:cell_methods = "time: mean" ;
		SNOBCMCL:_FillValue = 1.e+36f ;
		SNOBCMCL:missing_value = 1.e+36f ;
	float SNOBCMSL(time, lndgrid) ;
		SNOBCMSL:long_name = "mass of BC in top snow layer" ;
		SNOBCMSL:units = "kg/m2" ;
		SNOBCMSL:cell_methods = "time: mean" ;
		SNOBCMSL:_FillValue = 1.e+36f ;
		SNOBCMSL:missing_value = 1.e+36f ;
	float SNODSTMCL(time, lndgrid) ;
		SNODSTMCL:long_name = "mass of dust in snow column" ;
		SNODSTMCL:units = "kg/m2" ;
		SNODSTMCL:cell_methods = "time: mean" ;
		SNODSTMCL:_FillValue = 1.e+36f ;
		SNODSTMCL:missing_value = 1.e+36f ;
	float SNODSTMSL(time, lndgrid) ;
		SNODSTMSL:long_name = "mass of dust in top snow layer" ;
		SNODSTMSL:units = "kg/m2" ;
		SNODSTMSL:cell_methods = "time: mean" ;
		SNODSTMSL:_FillValue = 1.e+36f ;
		SNODSTMSL:missing_value = 1.e+36f ;
	float SNOINTABS(time, lndgrid) ;
		SNOINTABS:long_name = "Percent of incoming solar absorbed by lower snow layers" ;
		SNOINTABS:units = "%" ;
		SNOINTABS:cell_methods = "time: mean" ;
		SNOINTABS:_FillValue = 1.e+36f ;
		SNOINTABS:missing_value = 1.e+36f ;
	float SNOOCMCL(time, lndgrid) ;
		SNOOCMCL:long_name = "mass of OC in snow column" ;
		SNOOCMCL:units = "kg/m2" ;
		SNOOCMCL:cell_methods = "time: mean" ;
		SNOOCMCL:_FillValue = 1.e+36f ;
		SNOOCMCL:missing_value = 1.e+36f ;
	float SNOOCMSL(time, lndgrid) ;
		SNOOCMSL:long_name = "mass of OC in top snow layer" ;
		SNOOCMSL:units = "kg/m2" ;
		SNOOCMSL:cell_methods = "time: mean" ;
		SNOOCMSL:_FillValue = 1.e+36f ;
		SNOOCMSL:missing_value = 1.e+36f ;
	float SNOW(time, lndgrid) ;
		SNOW:long_name = "atmospheric snow" ;
		SNOW:units = "mm/s" ;
		SNOW:cell_methods = "time: mean" ;
		SNOW:_FillValue = 1.e+36f ;
		SNOW:missing_value = 1.e+36f ;
	float SNOWDP(time, lndgrid) ;
		SNOWDP:long_name = "gridcell mean snow height" ;
		SNOWDP:units = "m" ;
		SNOWDP:cell_methods = "time: mean" ;
		SNOWDP:_FillValue = 1.e+36f ;
		SNOWDP:missing_value = 1.e+36f ;
	float SNOWICE(time, lndgrid) ;
		SNOWICE:long_name = "snow ice" ;
		SNOWICE:units = "kg/m2" ;
		SNOWICE:cell_methods = "time: mean" ;
		SNOWICE:_FillValue = 1.e+36f ;
		SNOWICE:missing_value = 1.e+36f ;
	float SNOWLIQ(time, lndgrid) ;
		SNOWLIQ:long_name = "snow liquid water" ;
		SNOWLIQ:units = "kg/m2" ;
		SNOWLIQ:cell_methods = "time: mean" ;
		SNOWLIQ:_FillValue = 1.e+36f ;
		SNOWLIQ:missing_value = 1.e+36f ;
	float SNOW_DEPTH(time, lndgrid) ;
		SNOW_DEPTH:long_name = "snow height of snow covered area" ;
		SNOW_DEPTH:units = "m" ;
		SNOW_DEPTH:cell_methods = "time: mean" ;
		SNOW_DEPTH:_FillValue = 1.e+36f ;
		SNOW_DEPTH:missing_value = 1.e+36f ;
	float SNOW_SINKS(time, lndgrid) ;
		SNOW_SINKS:long_name = "snow sinks (liquid water)" ;
		SNOW_SINKS:units = "mm/s" ;
		SNOW_SINKS:cell_methods = "time: mean" ;
		SNOW_SINKS:_FillValue = 1.e+36f ;
		SNOW_SINKS:missing_value = 1.e+36f ;
	float SNOW_SOURCES(time, lndgrid) ;
		SNOW_SOURCES:long_name = "snow sources (liquid water)" ;
		SNOW_SOURCES:units = "mm/s" ;
		SNOW_SOURCES:cell_methods = "time: mean" ;
		SNOW_SOURCES:_FillValue = 1.e+36f ;
		SNOW_SOURCES:missing_value = 1.e+36f ;
	float SOIL1C(time, lndgrid) ;
		SOIL1C:long_name = "SOIL1 C" ;
		SOIL1C:units = "gC/m^2" ;
		SOIL1C:cell_methods = "time: mean" ;
		SOIL1C:_FillValue = 1.e+36f ;
		SOIL1C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL2C(time, lndgrid) ;
		SOIL1C_TO_SOIL2C:long_name = "decomp. of soil 1 C to soil 2 C" ;
		SOIL1C_TO_SOIL2C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL2C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL2C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL2C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL3C(time, lndgrid) ;
		SOIL1C_TO_SOIL3C:long_name = "decomp. of soil 1 C to soil 3 C" ;
		SOIL1C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL1C_vr(time, levdcmp, lndgrid) ;
		SOIL1C_vr:long_name = "SOIL1 C (vertically resolved)" ;
		SOIL1C_vr:units = "gC/m^3" ;
		SOIL1C_vr:cell_methods = "time: mean" ;
		SOIL1C_vr:_FillValue = 1.e+36f ;
		SOIL1C_vr:missing_value = 1.e+36f ;
	float SOIL1N(time, lndgrid) ;
		SOIL1N:long_name = "SOIL1 N" ;
		SOIL1N:units = "gN/m^2" ;
		SOIL1N:cell_methods = "time: mean" ;
		SOIL1N:_FillValue = 1.e+36f ;
		SOIL1N:missing_value = 1.e+36f ;
	float SOIL1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL1N_TNDNCY_VERT_TRANS:long_name = "soil 1 N tendency due to vertical transport" ;
		SOIL1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL2N(time, lndgrid) ;
		SOIL1N_TO_SOIL2N:long_name = "decomp. of soil 1 N to soil 2 N" ;
		SOIL1N_TO_SOIL2N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL2N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL2N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL2N:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL3N(time, lndgrid) ;
		SOIL1N_TO_SOIL3N:long_name = "decomp. of soil 1 N to soil 3 N" ;
		SOIL1N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL1N_vr(time, levdcmp, lndgrid) ;
		SOIL1N_vr:long_name = "SOIL1 N (vertically resolved)" ;
		SOIL1N_vr:units = "gN/m^3" ;
		SOIL1N_vr:cell_methods = "time: mean" ;
		SOIL1N_vr:_FillValue = 1.e+36f ;
		SOIL1N_vr:missing_value = 1.e+36f ;
	float SOIL1_HR_S2(time, lndgrid) ;
		SOIL1_HR_S2:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S2:units = "gC/m^2/s" ;
		SOIL1_HR_S2:cell_methods = "time: mean" ;
		SOIL1_HR_S2:_FillValue = 1.e+36f ;
		SOIL1_HR_S2:missing_value = 1.e+36f ;
	float SOIL1_HR_S3(time, lndgrid) ;
		SOIL1_HR_S3:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S3:units = "gC/m^2/s" ;
		SOIL1_HR_S3:cell_methods = "time: mean" ;
		SOIL1_HR_S3:_FillValue = 1.e+36f ;
		SOIL1_HR_S3:missing_value = 1.e+36f ;
	float SOIL2C(time, lndgrid) ;
		SOIL2C:long_name = "SOIL2 C" ;
		SOIL2C:units = "gC/m^2" ;
		SOIL2C:cell_methods = "time: mean" ;
		SOIL2C:_FillValue = 1.e+36f ;
		SOIL2C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL1C(time, lndgrid) ;
		SOIL2C_TO_SOIL1C:long_name = "decomp. of soil 2 C to soil 1 C" ;
		SOIL2C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL3C(time, lndgrid) ;
		SOIL2C_TO_SOIL3C:long_name = "decomp. of soil 2 C to soil 3 C" ;
		SOIL2C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL2C_vr(time, levdcmp, lndgrid) ;
		SOIL2C_vr:long_name = "SOIL2 C (vertically resolved)" ;
		SOIL2C_vr:units = "gC/m^3" ;
		SOIL2C_vr:cell_methods = "time: mean" ;
		SOIL2C_vr:_FillValue = 1.e+36f ;
		SOIL2C_vr:missing_value = 1.e+36f ;
	float SOIL2N(time, lndgrid) ;
		SOIL2N:long_name = "SOIL2 N" ;
		SOIL2N:units = "gN/m^2" ;
		SOIL2N:cell_methods = "time: mean" ;
		SOIL2N:_FillValue = 1.e+36f ;
		SOIL2N:missing_value = 1.e+36f ;
	float SOIL2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL2N_TNDNCY_VERT_TRANS:long_name = "soil 2 N tendency due to vertical transport" ;
		SOIL2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL1N(time, lndgrid) ;
		SOIL2N_TO_SOIL1N:long_name = "decomp. of soil 2 N to soil 1 N" ;
		SOIL2N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL3N(time, lndgrid) ;
		SOIL2N_TO_SOIL3N:long_name = "decomp. of soil 2 N to soil 3 N" ;
		SOIL2N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL2N_vr(time, levdcmp, lndgrid) ;
		SOIL2N_vr:long_name = "SOIL2 N (vertically resolved)" ;
		SOIL2N_vr:units = "gN/m^3" ;
		SOIL2N_vr:cell_methods = "time: mean" ;
		SOIL2N_vr:_FillValue = 1.e+36f ;
		SOIL2N_vr:missing_value = 1.e+36f ;
	float SOIL2_HR_S1(time, lndgrid) ;
		SOIL2_HR_S1:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S1:units = "gC/m^2/s" ;
		SOIL2_HR_S1:cell_methods = "time: mean" ;
		SOIL2_HR_S1:_FillValue = 1.e+36f ;
		SOIL2_HR_S1:missing_value = 1.e+36f ;
	float SOIL2_HR_S3(time, lndgrid) ;
		SOIL2_HR_S3:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S3:units = "gC/m^2/s" ;
		SOIL2_HR_S3:cell_methods = "time: mean" ;
		SOIL2_HR_S3:_FillValue = 1.e+36f ;
		SOIL2_HR_S3:missing_value = 1.e+36f ;
	float SOIL3C(time, lndgrid) ;
		SOIL3C:long_name = "SOIL3 C" ;
		SOIL3C:units = "gC/m^2" ;
		SOIL3C:cell_methods = "time: mean" ;
		SOIL3C:_FillValue = 1.e+36f ;
		SOIL3C:missing_value = 1.e+36f ;
	float SOIL3C_TO_SOIL1C(time, lndgrid) ;
		SOIL3C_TO_SOIL1C:long_name = "decomp. of soil 3 C to soil 1 C" ;
		SOIL3C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL3C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL3C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL3C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL3C_vr(time, levdcmp, lndgrid) ;
		SOIL3C_vr:long_name = "SOIL3 C (vertically resolved)" ;
		SOIL3C_vr:units = "gC/m^3" ;
		SOIL3C_vr:cell_methods = "time: mean" ;
		SOIL3C_vr:_FillValue = 1.e+36f ;
		SOIL3C_vr:missing_value = 1.e+36f ;
	float SOIL3N(time, lndgrid) ;
		SOIL3N:long_name = "SOIL3 N" ;
		SOIL3N:units = "gN/m^2" ;
		SOIL3N:cell_methods = "time: mean" ;
		SOIL3N:_FillValue = 1.e+36f ;
		SOIL3N:missing_value = 1.e+36f ;
	float SOIL3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL3N_TNDNCY_VERT_TRANS:long_name = "soil 3 N tendency due to vertical transport" ;
		SOIL3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL3N_TO_SOIL1N(time, lndgrid) ;
		SOIL3N_TO_SOIL1N:long_name = "decomp. of soil 3 N to soil 1 N" ;
		SOIL3N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL3N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL3N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL3N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL3N_vr(time, levdcmp, lndgrid) ;
		SOIL3N_vr:long_name = "SOIL3 N (vertically resolved)" ;
		SOIL3N_vr:units = "gN/m^3" ;
		SOIL3N_vr:cell_methods = "time: mean" ;
		SOIL3N_vr:_FillValue = 1.e+36f ;
		SOIL3N_vr:missing_value = 1.e+36f ;
	float SOIL3_HR(time, lndgrid) ;
		SOIL3_HR:long_name = "Het. Resp. from soil 3" ;
		SOIL3_HR:units = "gC/m^2/s" ;
		SOIL3_HR:cell_methods = "time: mean" ;
		SOIL3_HR:_FillValue = 1.e+36f ;
		SOIL3_HR:missing_value = 1.e+36f ;
	float SOILC(time, lndgrid) ;
		SOILC:long_name = "soil C" ;
		SOILC:units = "gC/m^2" ;
		SOILC:cell_methods = "time: mean" ;
		SOILC:_FillValue = 1.e+36f ;
		SOILC:missing_value = 1.e+36f ;
	float SOILC_HR(time, lndgrid) ;
		SOILC_HR:long_name = "soil C heterotrophic respiration" ;
		SOILC_HR:units = "gC/m^2/s" ;
		SOILC_HR:cell_methods = "time: mean" ;
		SOILC_HR:_FillValue = 1.e+36f ;
		SOILC_HR:missing_value = 1.e+36f ;
	float SOILC_LOSS(time, lndgrid) ;
		SOILC_LOSS:long_name = "soil C loss" ;
		SOILC_LOSS:units = "gC/m^2/s" ;
		SOILC_LOSS:cell_methods = "time: mean" ;
		SOILC_LOSS:_FillValue = 1.e+36f ;
		SOILC_LOSS:missing_value = 1.e+36f ;
	float SOILICE(time, levgrnd, lndgrid) ;
		SOILICE:long_name = "soil ice (vegetated landunits only)" ;
		SOILICE:units = "kg/m2" ;
		SOILICE:cell_methods = "time: mean" ;
		SOILICE:_FillValue = 1.e+36f ;
		SOILICE:missing_value = 1.e+36f ;
	float SOILLIQ(time, levgrnd, lndgrid) ;
		SOILLIQ:long_name = "soil liquid water (vegetated landunits only)" ;
		SOILLIQ:units = "kg/m2" ;
		SOILLIQ:cell_methods = "time: mean" ;
		SOILLIQ:_FillValue = 1.e+36f ;
		SOILLIQ:missing_value = 1.e+36f ;
	float SOILPSI(time, levgrnd, lndgrid) ;
		SOILPSI:long_name = "soil water potential in each soil layer" ;
		SOILPSI:units = "MPa" ;
		SOILPSI:cell_methods = "time: mean" ;
		SOILPSI:_FillValue = 1.e+36f ;
		SOILPSI:missing_value = 1.e+36f ;
	float SOILWATER_10CM(time, lndgrid) ;
		SOILWATER_10CM:long_name = "soil liquid water + ice in top 10cm of soil (veg landunits only)" ;
		SOILWATER_10CM:units = "kg/m2" ;
		SOILWATER_10CM:cell_methods = "time: mean" ;
		SOILWATER_10CM:_FillValue = 1.e+36f ;
		SOILWATER_10CM:missing_value = 1.e+36f ;
	float SOMC_FIRE(time, lndgrid) ;
		SOMC_FIRE:long_name = "C loss due to peat burning" ;
		SOMC_FIRE:units = "gC/m^2/s" ;
		SOMC_FIRE:cell_methods = "time: mean" ;
		SOMC_FIRE:_FillValue = 1.e+36f ;
		SOMC_FIRE:missing_value = 1.e+36f ;
	float SOMHR(time, lndgrid) ;
		SOMHR:long_name = "soil organic matter heterotrophic respiration" ;
		SOMHR:units = "gC/m^2/s" ;
		SOMHR:cell_methods = "time: mean" ;
		SOMHR:_FillValue = 1.e+36f ;
		SOMHR:missing_value = 1.e+36f ;
	float SOM_C_LEACHED(time, lndgrid) ;
		SOM_C_LEACHED:long_name = "total flux of C from SOM pools due to leaching" ;
		SOM_C_LEACHED:units = "gC/m^2/s" ;
		SOM_C_LEACHED:cell_methods = "time: mean" ;
		SOM_C_LEACHED:_FillValue = 1.e+36f ;
		SOM_C_LEACHED:missing_value = 1.e+36f ;
	float SR(time, lndgrid) ;
		SR:long_name = "total soil respiration (HR + root resp)" ;
		SR:units = "gC/m^2/s" ;
		SR:cell_methods = "time: mean" ;
		SR:_FillValue = 1.e+36f ;
		SR:missing_value = 1.e+36f ;
	float STORVEGC(time, lndgrid) ;
		STORVEGC:long_name = "stored vegetation carbon, excluding cpool" ;
		STORVEGC:units = "gC/m^2" ;
		STORVEGC:cell_methods = "time: mean" ;
		STORVEGC:_FillValue = 1.e+36f ;
		STORVEGC:missing_value = 1.e+36f ;
	float STORVEGN(time, lndgrid) ;
		STORVEGN:long_name = "stored vegetation nitrogen" ;
		STORVEGN:units = "gN/m^2" ;
		STORVEGN:cell_methods = "time: mean" ;
		STORVEGN:_FillValue = 1.e+36f ;
		STORVEGN:missing_value = 1.e+36f ;
	float SUPPLEMENT_TO_SMINN(time, lndgrid) ;
		SUPPLEMENT_TO_SMINN:long_name = "supplemental N supply" ;
		SUPPLEMENT_TO_SMINN:units = "gN/m^2/s" ;
		SUPPLEMENT_TO_SMINN:cell_methods = "time: mean" ;
		SUPPLEMENT_TO_SMINN:_FillValue = 1.e+36f ;
		SUPPLEMENT_TO_SMINN:missing_value = 1.e+36f ;
	float SoilAlpha(time, lndgrid) ;
		SoilAlpha:long_name = "factor limiting ground evap" ;
		SoilAlpha:units = "unitless" ;
		SoilAlpha:cell_methods = "time: mean" ;
		SoilAlpha:_FillValue = 1.e+36f ;
		SoilAlpha:missing_value = 1.e+36f ;
	float SoilAlpha_U(time, lndgrid) ;
		SoilAlpha_U:long_name = "urban factor limiting ground evap" ;
		SoilAlpha_U:units = "unitless" ;
		SoilAlpha_U:cell_methods = "time: mean" ;
		SoilAlpha_U:_FillValue = 1.e+36f ;
		SoilAlpha_U:missing_value = 1.e+36f ;
	float TAUX(time, lndgrid) ;
		TAUX:long_name = "zonal surface stress" ;
		TAUX:units = "kg/m/s^2" ;
		TAUX:cell_methods = "time: mean" ;
		TAUX:_FillValue = 1.e+36f ;
		TAUX:missing_value = 1.e+36f ;
	float TAUY(time, lndgrid) ;
		TAUY:long_name = "meridional surface stress" ;
		TAUY:units = "kg/m/s^2" ;
		TAUY:cell_methods = "time: mean" ;
		TAUY:_FillValue = 1.e+36f ;
		TAUY:missing_value = 1.e+36f ;
	float TBOT(time, lndgrid) ;
		TBOT:long_name = "atmospheric air temperature" ;
		TBOT:units = "K" ;
		TBOT:cell_methods = "time: mean" ;
		TBOT:_FillValue = 1.e+36f ;
		TBOT:missing_value = 1.e+36f ;
	float TBUILD(time, lndgrid) ;
		TBUILD:long_name = "internal urban building temperature" ;
		TBUILD:units = "K" ;
		TBUILD:cell_methods = "time: mean" ;
		TBUILD:_FillValue = 1.e+36f ;
		TBUILD:missing_value = 1.e+36f ;
	float TG(time, lndgrid) ;
		TG:long_name = "ground temperature" ;
		TG:units = "K" ;
		TG:cell_methods = "time: mean" ;
		TG:_FillValue = 1.e+36f ;
		TG:missing_value = 1.e+36f ;
	float TG_R(time, lndgrid) ;
		TG_R:long_name = "Rural ground temperature" ;
		TG_R:units = "K" ;
		TG_R:cell_methods = "time: mean" ;
		TG_R:_FillValue = 1.e+36f ;
		TG_R:missing_value = 1.e+36f ;
	float TG_U(time, lndgrid) ;
		TG_U:long_name = "Urban ground temperature" ;
		TG_U:units = "K" ;
		TG_U:cell_methods = "time: mean" ;
		TG_U:_FillValue = 1.e+36f ;
		TG_U:missing_value = 1.e+36f ;
	float TH2OSFC(time, lndgrid) ;
		TH2OSFC:long_name = "surface water temperature" ;
		TH2OSFC:units = "K" ;
		TH2OSFC:cell_methods = "time: mean" ;
		TH2OSFC:_FillValue = 1.e+36f ;
		TH2OSFC:missing_value = 1.e+36f ;
	float THBOT(time, lndgrid) ;
		THBOT:long_name = "atmospheric air potential temperature" ;
		THBOT:units = "K" ;
		THBOT:cell_methods = "time: mean" ;
		THBOT:_FillValue = 1.e+36f ;
		THBOT:missing_value = 1.e+36f ;
	float TKE1(time, lndgrid) ;
		TKE1:long_name = "top lake level eddy thermal conductivity" ;
		TKE1:units = "W/(mK)" ;
		TKE1:cell_methods = "time: mean" ;
		TKE1:_FillValue = 1.e+36f ;
		TKE1:missing_value = 1.e+36f ;
	float TLAI(time, lndgrid) ;
		TLAI:long_name = "total projected leaf area index" ;
		TLAI:units = "none" ;
		TLAI:cell_methods = "time: mean" ;
		TLAI:_FillValue = 1.e+36f ;
		TLAI:missing_value = 1.e+36f ;
	float TLAKE(time, levlak, lndgrid) ;
		TLAKE:long_name = "lake temperature" ;
		TLAKE:units = "K" ;
		TLAKE:cell_methods = "time: mean" ;
		TLAKE:_FillValue = 1.e+36f ;
		TLAKE:missing_value = 1.e+36f ;
	float TOTCOLC(time, lndgrid) ;
		TOTCOLC:long_name = "total column carbon, incl veg and cpool" ;
		TOTCOLC:units = "gC/m^2" ;
		TOTCOLC:cell_methods = "time: mean" ;
		TOTCOLC:_FillValue = 1.e+36f ;
		TOTCOLC:missing_value = 1.e+36f ;
	float TOTCOLCH4(time, lndgrid) ;
		TOTCOLCH4:long_name = "total belowground CH4, (0 for non-lake special landunits)" ;
		TOTCOLCH4:units = "gC/m2" ;
		TOTCOLCH4:cell_methods = "time: mean" ;
		TOTCOLCH4:_FillValue = 1.e+36f ;
		TOTCOLCH4:missing_value = 1.e+36f ;
	float TOTCOLN(time, lndgrid) ;
		TOTCOLN:long_name = "total column-level N" ;
		TOTCOLN:units = "gN/m^2" ;
		TOTCOLN:cell_methods = "time: mean" ;
		TOTCOLN:_FillValue = 1.e+36f ;
		TOTCOLN:missing_value = 1.e+36f ;
	float TOTECOSYSC(time, lndgrid) ;
		TOTECOSYSC:long_name = "total ecosystem carbon, incl veg but excl cpool" ;
		TOTECOSYSC:units = "gC/m^2" ;
		TOTECOSYSC:cell_methods = "time: mean" ;
		TOTECOSYSC:_FillValue = 1.e+36f ;
		TOTECOSYSC:missing_value = 1.e+36f ;
	float TOTECOSYSN(time, lndgrid) ;
		TOTECOSYSN:long_name = "total ecosystem N" ;
		TOTECOSYSN:units = "gN/m^2" ;
		TOTECOSYSN:cell_methods = "time: mean" ;
		TOTECOSYSN:_FillValue = 1.e+36f ;
		TOTECOSYSN:missing_value = 1.e+36f ;
	float TOTLITC(time, lndgrid) ;
		TOTLITC:long_name = "total litter carbon" ;
		TOTLITC:units = "gC/m^2" ;
		TOTLITC:cell_methods = "time: mean" ;
		TOTLITC:_FillValue = 1.e+36f ;
		TOTLITC:missing_value = 1.e+36f ;
	float TOTLITC_1m(time, lndgrid) ;
		TOTLITC_1m:long_name = "total litter carbon to 1 meter depth" ;
		TOTLITC_1m:units = "gC/m^2" ;
		TOTLITC_1m:cell_methods = "time: mean" ;
		TOTLITC_1m:_FillValue = 1.e+36f ;
		TOTLITC_1m:missing_value = 1.e+36f ;
	float TOTLITN(time, lndgrid) ;
		TOTLITN:long_name = "total litter N" ;
		TOTLITN:units = "gN/m^2" ;
		TOTLITN:cell_methods = "time: mean" ;
		TOTLITN:_FillValue = 1.e+36f ;
		TOTLITN:missing_value = 1.e+36f ;
	float TOTLITN_1m(time, lndgrid) ;
		TOTLITN_1m:long_name = "total litter N to 1 meter" ;
		TOTLITN_1m:units = "gN/m^2" ;
		TOTLITN_1m:cell_methods = "time: mean" ;
		TOTLITN_1m:_FillValue = 1.e+36f ;
		TOTLITN_1m:missing_value = 1.e+36f ;
	float TOTPFTC(time, lndgrid) ;
		TOTPFTC:long_name = "total pft-level carbon, including cpool" ;
		TOTPFTC:units = "gC/m^2" ;
		TOTPFTC:cell_methods = "time: mean" ;
		TOTPFTC:_FillValue = 1.e+36f ;
		TOTPFTC:missing_value = 1.e+36f ;
	float TOTPFTN(time, lndgrid) ;
		TOTPFTN:long_name = "total PFT-level nitrogen" ;
		TOTPFTN:units = "gN/m^2" ;
		TOTPFTN:cell_methods = "time: mean" ;
		TOTPFTN:_FillValue = 1.e+36f ;
		TOTPFTN:missing_value = 1.e+36f ;
	float TOTPRODC(time, lndgrid) ;
		TOTPRODC:long_name = "total wood product C" ;
		TOTPRODC:units = "gC/m^2" ;
		TOTPRODC:cell_methods = "time: mean" ;
		TOTPRODC:_FillValue = 1.e+36f ;
		TOTPRODC:missing_value = 1.e+36f ;
	float TOTPRODN(time, lndgrid) ;
		TOTPRODN:long_name = "total wood product N" ;
		TOTPRODN:units = "gN/m^2" ;
		TOTPRODN:cell_methods = "time: mean" ;
		TOTPRODN:_FillValue = 1.e+36f ;
		TOTPRODN:missing_value = 1.e+36f ;
	float TOTSOMC(time, lndgrid) ;
		TOTSOMC:long_name = "total soil organic matter carbon" ;
		TOTSOMC:units = "gC/m^2" ;
		TOTSOMC:cell_methods = "time: mean" ;
		TOTSOMC:_FillValue = 1.e+36f ;
		TOTSOMC:missing_value = 1.e+36f ;
	float TOTSOMC_1m(time, lndgrid) ;
		TOTSOMC_1m:long_name = "total soil organic matter carbon to 1 meter depth" ;
		TOTSOMC_1m:units = "gC/m^2" ;
		TOTSOMC_1m:cell_methods = "time: mean" ;
		TOTSOMC_1m:_FillValue = 1.e+36f ;
		TOTSOMC_1m:missing_value = 1.e+36f ;
	float TOTSOMN(time, lndgrid) ;
		TOTSOMN:long_name = "total soil organic matter N" ;
		TOTSOMN:units = "gN/m^2" ;
		TOTSOMN:cell_methods = "time: mean" ;
		TOTSOMN:_FillValue = 1.e+36f ;
		TOTSOMN:missing_value = 1.e+36f ;
	float TOTSOMN_1m(time, lndgrid) ;
		TOTSOMN_1m:long_name = "total soil organic matter N to 1 meter" ;
		TOTSOMN_1m:units = "gN/m^2" ;
		TOTSOMN_1m:cell_methods = "time: mean" ;
		TOTSOMN_1m:_FillValue = 1.e+36f ;
		TOTSOMN_1m:missing_value = 1.e+36f ;
	float TOTVEGC(time, lndgrid) ;
		TOTVEGC:long_name = "total vegetation carbon, excluding cpool" ;
		TOTVEGC:units = "gC/m^2" ;
		TOTVEGC:cell_methods = "time: mean" ;
		TOTVEGC:_FillValue = 1.e+36f ;
		TOTVEGC:missing_value = 1.e+36f ;
	float TOTVEGN(time, lndgrid) ;
		TOTVEGN:long_name = "total vegetation nitrogen" ;
		TOTVEGN:units = "gN/m^2" ;
		TOTVEGN:cell_methods = "time: mean" ;
		TOTVEGN:_FillValue = 1.e+36f ;
		TOTVEGN:missing_value = 1.e+36f ;
	float TREFMNAV(time, lndgrid) ;
		TREFMNAV:long_name = "daily minimum of average 2-m temperature" ;
		TREFMNAV:units = "K" ;
		TREFMNAV:cell_methods = "time: mean" ;
		TREFMNAV:_FillValue = 1.e+36f ;
		TREFMNAV:missing_value = 1.e+36f ;
	float TREFMNAV_R(time, lndgrid) ;
		TREFMNAV_R:long_name = "Rural daily minimum of average 2-m temperature" ;
		TREFMNAV_R:units = "K" ;
		TREFMNAV_R:cell_methods = "time: mean" ;
		TREFMNAV_R:_FillValue = 1.e+36f ;
		TREFMNAV_R:missing_value = 1.e+36f ;
	float TREFMNAV_U(time, lndgrid) ;
		TREFMNAV_U:long_name = "Urban daily minimum of average 2-m temperature" ;
		TREFMNAV_U:units = "K" ;
		TREFMNAV_U:cell_methods = "time: mean" ;
		TREFMNAV_U:_FillValue = 1.e+36f ;
		TREFMNAV_U:missing_value = 1.e+36f ;
	float TREFMXAV(time, lndgrid) ;
		TREFMXAV:long_name = "daily maximum of average 2-m temperature" ;
		TREFMXAV:units = "K" ;
		TREFMXAV:cell_methods = "time: mean" ;
		TREFMXAV:_FillValue = 1.e+36f ;
		TREFMXAV:missing_value = 1.e+36f ;
	float TREFMXAV_R(time, lndgrid) ;
		TREFMXAV_R:long_name = "Rural daily maximum of average 2-m temperature" ;
		TREFMXAV_R:units = "K" ;
		TREFMXAV_R:cell_methods = "time: mean" ;
		TREFMXAV_R:_FillValue = 1.e+36f ;
		TREFMXAV_R:missing_value = 1.e+36f ;
	float TREFMXAV_U(time, lndgrid) ;
		TREFMXAV_U:long_name = "Urban daily maximum of average 2-m temperature" ;
		TREFMXAV_U:units = "K" ;
		TREFMXAV_U:cell_methods = "time: mean" ;
		TREFMXAV_U:_FillValue = 1.e+36f ;
		TREFMXAV_U:missing_value = 1.e+36f ;
	float TSA(time, lndgrid) ;
		TSA:long_name = "2m air temperature" ;
		TSA:units = "K" ;
		TSA:cell_methods = "time: mean" ;
		TSA:_FillValue = 1.e+36f ;
		TSA:missing_value = 1.e+36f ;
	float TSAI(time, lndgrid) ;
		TSAI:long_name = "total projected stem area index" ;
		TSAI:units = "none" ;
		TSAI:cell_methods = "time: mean" ;
		TSAI:_FillValue = 1.e+36f ;
		TSAI:missing_value = 1.e+36f ;
	float TSA_R(time, lndgrid) ;
		TSA_R:long_name = "Rural 2m air temperature" ;
		TSA_R:units = "K" ;
		TSA_R:cell_methods = "time: mean" ;
		TSA_R:_FillValue = 1.e+36f ;
		TSA_R:missing_value = 1.e+36f ;
	float TSA_U(time, lndgrid) ;
		TSA_U:long_name = "Urban 2m air temperature" ;
		TSA_U:units = "K" ;
		TSA_U:cell_methods = "time: mean" ;
		TSA_U:_FillValue = 1.e+36f ;
		TSA_U:missing_value = 1.e+36f ;
	float TSOI(time, levgrnd, lndgrid) ;
		TSOI:long_name = "soil temperature (vegetated landunits only)" ;
		TSOI:units = "K" ;
		TSOI:cell_methods = "time: mean" ;
		TSOI:_FillValue = 1.e+36f ;
		TSOI:missing_value = 1.e+36f ;
	float TSOI_10CM(time, lndgrid) ;
		TSOI_10CM:long_name = "soil temperature in top 10cm of soil" ;
		TSOI_10CM:units = "K" ;
		TSOI_10CM:cell_methods = "time: mean" ;
		TSOI_10CM:_FillValue = 1.e+36f ;
		TSOI_10CM:missing_value = 1.e+36f ;
	float TSOI_ICE(time, levgrnd, lndgrid) ;
		TSOI_ICE:long_name = "soil temperature (ice landunits only)" ;
		TSOI_ICE:units = "K" ;
		TSOI_ICE:cell_methods = "time: mean" ;
		TSOI_ICE:_FillValue = 1.e+36f ;
		TSOI_ICE:missing_value = 1.e+36f ;
	float TV(time, lndgrid) ;
		TV:long_name = "vegetation temperature" ;
		TV:units = "K" ;
		TV:cell_methods = "time: mean" ;
		TV:_FillValue = 1.e+36f ;
		TV:missing_value = 1.e+36f ;
	float TWS(time, lndgrid) ;
		TWS:long_name = "total water storage" ;
		TWS:units = "mm" ;
		TWS:cell_methods = "time: mean" ;
		TWS:_FillValue = 1.e+36f ;
		TWS:missing_value = 1.e+36f ;
	float T_SCALAR(time, levdcmp, lndgrid) ;
		T_SCALAR:long_name = "temperature inhibition of decomposition" ;
		T_SCALAR:units = "unitless" ;
		T_SCALAR:cell_methods = "time: mean" ;
		T_SCALAR:_FillValue = 1.e+36f ;
		T_SCALAR:missing_value = 1.e+36f ;
	float U10(time, lndgrid) ;
		U10:long_name = "10-m wind" ;
		U10:units = "m/s" ;
		U10:cell_methods = "time: mean" ;
		U10:_FillValue = 1.e+36f ;
		U10:missing_value = 1.e+36f ;
	float URBAN_AC(time, lndgrid) ;
		URBAN_AC:long_name = "urban air conditioning flux" ;
		URBAN_AC:units = "W/m^2" ;
		URBAN_AC:cell_methods = "time: mean" ;
		URBAN_AC:_FillValue = 1.e+36f ;
		URBAN_AC:missing_value = 1.e+36f ;
	float URBAN_HEAT(time, lndgrid) ;
		URBAN_HEAT:long_name = "urban heating flux" ;
		URBAN_HEAT:units = "W/m^2" ;
		URBAN_HEAT:cell_methods = "time: mean" ;
		URBAN_HEAT:_FillValue = 1.e+36f ;
		URBAN_HEAT:missing_value = 1.e+36f ;
	float VOCFLXT(time, lndgrid) ;
		VOCFLXT:long_name = "total VOC flux into atmosphere" ;
		VOCFLXT:units = "moles/m2/sec" ;
		VOCFLXT:cell_methods = "time: mean" ;
		VOCFLXT:_FillValue = 1.e+36f ;
		VOCFLXT:missing_value = 1.e+36f ;
	float VOLR(time, lndgrid) ;
		VOLR:long_name = "river channel water storage" ;
		VOLR:units = "m3" ;
		VOLR:cell_methods = "time: mean" ;
		VOLR:_FillValue = 1.e+36f ;
		VOLR:missing_value = 1.e+36f ;
	float WA(time, lndgrid) ;
		WA:long_name = "water in the unconfined aquifer (vegetated landunits only)" ;
		WA:units = "mm" ;
		WA:cell_methods = "time: mean" ;
		WA:_FillValue = 1.e+36f ;
		WA:missing_value = 1.e+36f ;
	float WASTEHEAT(time, lndgrid) ;
		WASTEHEAT:long_name = "sensible heat flux from heating/cooling sources of urban waste heat" ;
		WASTEHEAT:units = "W/m^2" ;
		WASTEHEAT:cell_methods = "time: mean" ;
		WASTEHEAT:_FillValue = 1.e+36f ;
		WASTEHEAT:missing_value = 1.e+36f ;
	float WF(time, lndgrid) ;
		WF:long_name = "soil water as frac. of whc for top 0.05 m" ;
		WF:units = "proportion" ;
		WF:cell_methods = "time: mean" ;
		WF:_FillValue = 1.e+36f ;
		WF:missing_value = 1.e+36f ;
	float WIND(time, lndgrid) ;
		WIND:long_name = "atmospheric wind velocity magnitude" ;
		WIND:units = "m/s" ;
		WIND:cell_methods = "time: mean" ;
		WIND:_FillValue = 1.e+36f ;
		WIND:missing_value = 1.e+36f ;
	float WOODC(time, lndgrid) ;
		WOODC:long_name = "wood C" ;
		WOODC:units = "gC/m^2" ;
		WOODC:cell_methods = "time: mean" ;
		WOODC:_FillValue = 1.e+36f ;
		WOODC:missing_value = 1.e+36f ;
	float WOODC_ALLOC(time, lndgrid) ;
		WOODC_ALLOC:long_name = "wood C allocation" ;
		WOODC_ALLOC:units = "gC/m^2/s" ;
		WOODC_ALLOC:cell_methods = "time: mean" ;
		WOODC_ALLOC:_FillValue = 1.e+36f ;
		WOODC_ALLOC:missing_value = 1.e+36f ;
	float WOODC_LOSS(time, lndgrid) ;
		WOODC_LOSS:long_name = "wood C loss" ;
		WOODC_LOSS:units = "gC/m^2/s" ;
		WOODC_LOSS:cell_methods = "time: mean" ;
		WOODC_LOSS:_FillValue = 1.e+36f ;
		WOODC_LOSS:missing_value = 1.e+36f ;
	float WOOD_HARVESTC(time, lndgrid) ;
		WOOD_HARVESTC:long_name = "wood harvest carbon (to product pools)" ;
		WOOD_HARVESTC:units = "gC/m^2/s" ;
		WOOD_HARVESTC:cell_methods = "time: mean" ;
		WOOD_HARVESTC:_FillValue = 1.e+36f ;
		WOOD_HARVESTC:missing_value = 1.e+36f ;
	float WOOD_HARVESTN(time, lndgrid) ;
		WOOD_HARVESTN:long_name = "wood harvest N (to product pools)" ;
		WOOD_HARVESTN:units = "gN/m^2/s" ;
		WOOD_HARVESTN:cell_methods = "time: mean" ;
		WOOD_HARVESTN:_FillValue = 1.e+36f ;
		WOOD_HARVESTN:missing_value = 1.e+36f ;
	float WTGQ(time, lndgrid) ;
		WTGQ:long_name = "surface tracer conductance" ;
		WTGQ:units = "m/s" ;
		WTGQ:cell_methods = "time: mean" ;
		WTGQ:_FillValue = 1.e+36f ;
		WTGQ:missing_value = 1.e+36f ;
	float W_SCALAR(time, levdcmp, lndgrid) ;
		W_SCALAR:long_name = "Moisture (dryness) inhibition of decomposition" ;
		W_SCALAR:units = "unitless" ;
		W_SCALAR:cell_methods = "time: mean" ;
		W_SCALAR:_FillValue = 1.e+36f ;
		W_SCALAR:missing_value = 1.e+36f ;
	float XSMRPOOL(time, lndgrid) ;
		XSMRPOOL:long_name = "temporary photosynthate C pool" ;
		XSMRPOOL:units = "gC/m^2" ;
		XSMRPOOL:cell_methods = "time: mean" ;
		XSMRPOOL:_FillValue = 1.e+36f ;
		XSMRPOOL:missing_value = 1.e+36f ;
	float XSMRPOOL_RECOVER(time, lndgrid) ;
		XSMRPOOL_RECOVER:long_name = "C flux assigned to recovery of negative xsmrpool" ;
		XSMRPOOL_RECOVER:units = "gC/m^2/s" ;
		XSMRPOOL_RECOVER:cell_methods = "time: mean" ;
		XSMRPOOL_RECOVER:_FillValue = 1.e+36f ;
		XSMRPOOL_RECOVER:missing_value = 1.e+36f ;
	float ZBOT(time, lndgrid) ;
		ZBOT:long_name = "atmospheric reference height" ;
		ZBOT:units = "m" ;
		ZBOT:cell_methods = "time: mean" ;
		ZBOT:_FillValue = 1.e+36f ;
		ZBOT:missing_value = 1.e+36f ;
	float ZWT(time, lndgrid) ;
		ZWT:long_name = "water table depth (vegetated landunits only)" ;
		ZWT:units = "m" ;
		ZWT:cell_methods = "time: mean" ;
		ZWT:_FillValue = 1.e+36f ;
		ZWT:missing_value = 1.e+36f ;
	float ZWT_CH4_UNSAT(time, lndgrid) ;
		ZWT_CH4_UNSAT:long_name = "depth of water table for methane production used in non-inundated area" ;
		ZWT_CH4_UNSAT:units = "m" ;
		ZWT_CH4_UNSAT:cell_methods = "time: mean" ;
		ZWT_CH4_UNSAT:_FillValue = 1.e+36f ;
		ZWT_CH4_UNSAT:missing_value = 1.e+36f ;
	float ZWT_PERCH(time, lndgrid) ;
		ZWT_PERCH:long_name = "perched water table depth (vegetated landunits only)" ;
		ZWT_PERCH:units = "m" ;
		ZWT_PERCH:cell_methods = "time: mean" ;
		ZWT_PERCH:_FillValue = 1.e+36f ;
		ZWT_PERCH:missing_value = 1.e+36f ;
	float o2_decomp_depth_unsat(time, levgrnd, lndgrid) ;
		o2_decomp_depth_unsat:long_name = "o2_decomp_depth_unsat" ;
		o2_decomp_depth_unsat:units = "mol/m3/2" ;
		o2_decomp_depth_unsat:cell_methods = "time: mean" ;
		o2_decomp_depth_unsat:_FillValue = 1.e+36f ;
		o2_decomp_depth_unsat:missing_value = 1.e+36f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "created on 08/20/14 15:53:41" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "userdefined" ;
		:username = "gbisht" ;
		:version = "" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "ugrid-13x26x10-surface-subsurface-th-noice-dec-NGEE_SiteB" ;
		:Surface_dataset = "surfdata_13x26pt_US-Brw_simyr1850.nc" ;
		:Initial_conditions_dataset = "arbitrary initialization" ;
		:PFT_physiological_constants_dataset = "clm_params.c140423.nc" ;
		:ltype_vegetated_or_bare_soil = 1 ;
		:ltype_crop = 2 ;
		:ltype_landice = 3 ;
		:ltype_landice_multiple_elevation_classes = 4 ;
		:ltype_deep_lake = 5 ;
		:ltype_wetland = 6 ;
		:ltype_urban_tbd = 7 ;
		:ltype_urban_hd = 8 ;
		:ltype_urban_md = 9 ;
		:natpft_not_vegetated = 1 ;
		:natpft_needleleaf_evergreen_temperate_tree = 2 ;
		:natpft_needleleaf_evergreen_boreal_tree = 3 ;
		:natpft_needleleaf_deciduous_boreal_tree = 4 ;
		:natpft_broadleaf_evergreen_tropical_tree = 5 ;
		:natpft_broadleaf_evergreen_temperate_tree = 6 ;
		:natpft_broadleaf_deciduous_tropical_tree = 7 ;
		:natpft_broadleaf_deciduous_temperate_tree = 8 ;
		:natpft_broadleaf_deciduous_boreal_tree = 9 ;
		:natpft_broadleaf_evergreen_shrub = 10 ;
		:natpft_broadleaf_deciduous_temperate_shrub = 11 ;
		:natpft_broadleaf_deciduous_boreal_shrub = 12 ;
		:natpft_c3_arctic_grass = 13 ;
		:natpft_c3_non-arctic_grass = 14 ;
		:natpft_c4_grass = 15 ;
		:natpft_c3_crop = 16 ;
		:natpft_c3_irrigated = 17 ;
		:Time_constant_3Dvars_filename = "./ugrid-13x26x10-surface-subsurface-th-noice-dec-NGEE_SiteB.clm2.h0.0001-01-01-00000.nc" ;
		:Time_constant_3Dvars = "ZSOI:DZSOI:WATSAT:SUCSAT:BSW:HKSAT:ZLAKE:DZLAKE" ;
data:

 levgrnd = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 levlak = 0.05, 0.6, 2.1, 4.6, 8.1, 12.6, 18.6, 25.6, 34.325, 44.775 ;

 levdcmp = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 time = 1 ;

 mcdate = 10102 ;

 mcsec = 0 ;

 mdcur = 1 ;

 mscur = 0 ;

 nstep = 48 ;

 time_bounds =
  0, 1 ;

 date_written =
  "08/20/14" ;

 time_written =
  "15:53:41" ;

 lon = -156.6089, -156.6089, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6083, -156.6082, -156.608, -156.608, -156.6078, -156.6078, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, 
    -156.6069, -156.6069, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6063, -156.6062, -156.6089, -156.6089, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6083, -156.6082, -156.608, -156.608, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6074, -156.6073, 
    -156.6071, -156.6071, -156.6069, -156.6069, -156.6067, -156.6066, 
    -156.6065, -156.6064, -156.6063, -156.6062, -156.6089, -156.6089, 
    -156.6087, -156.6086, -156.6085, -156.6084, -156.6083, -156.6082, 
    -156.608, -156.608, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6074, -156.6073, -156.6071, -156.6071, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6065, -156.6064, -156.6062, -156.6062, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6082, -156.6082, -156.608, -156.608, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6071, -156.6071, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6062, -156.6062, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6082, -156.6082, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6073, -156.6073, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6067, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6062, -156.6089, -156.6088, 
    -156.6087, -156.6086, -156.6084, -156.6084, -156.6082, -156.6082, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6073, -156.6073, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6064, -156.6064, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6084, -156.6084, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6073, -156.6073, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6064, -156.6064, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6084, -156.6084, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6075, -156.6075, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6061, -156.6089, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6084, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6075, -156.6075, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6066, -156.6066, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6086, -156.6086, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6075, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6066, -156.6066, -156.6064, -156.6063, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6086, -156.6086, 
    -156.6084, -156.6083, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6077, -156.6077, -156.6075, -156.6074, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6068, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6063, -156.6062, -156.6061, -156.6088, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6083, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6077, -156.6077, -156.6075, -156.6074, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6068, -156.6068, 
    -156.6066, -156.6065, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6088, -156.6088, -156.6086, -156.6085, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.6079, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6068, -156.6068, -156.6066, -156.6065, -156.6064, -156.6063, 
    -156.6062, -156.6061 ;

 lat = 71.27904, 71.27901, 71.27903, 71.27901, 71.27901, 71.27903, 71.27901, 
    71.27903, 71.279, 71.27902, 71.27902, 71.279, 71.27899, 71.27901, 
    71.27901, 71.27899, 71.27899, 71.27901, 71.27898, 71.27901, 71.27901, 
    71.27898, 71.27901, 71.27898, 71.27898, 71.279, 71.27911, 71.27908, 
    71.27911, 71.27908, 71.27908, 71.2791, 71.27908, 71.2791, 71.2791, 
    71.27907, 71.27907, 71.27909, 71.27909, 71.27907, 71.27909, 71.27906, 
    71.27906, 71.27908, 71.27906, 71.27908, 71.27905, 71.27908, 71.27908, 
    71.27905, 71.27908, 71.27905, 71.27915, 71.27918, 71.27915, 71.27917, 
    71.27917, 71.27915, 71.27917, 71.27914, 71.27914, 71.27917, 71.27914, 
    71.27917, 71.27916, 71.27914, 71.27914, 71.27916, 71.27914, 71.27916, 
    71.27913, 71.27915, 71.27913, 71.27915, 71.27915, 71.27912, 71.27914, 
    71.27912, 71.27923, 71.27925, 71.27923, 71.27925, 71.27924, 71.27922, 
    71.27922, 71.27924, 71.27921, 71.27924, 71.27921, 71.27924, 71.27924, 
    71.27921, 71.27921, 71.27923, 71.27923, 71.27921, 71.27923, 71.2792, 
    71.27922, 71.2792, 71.27922, 71.2792, 71.27922, 71.27919, 71.27932, 
    71.2793, 71.2793, 71.27932, 71.2793, 71.27932, 71.27931, 71.27929, 
    71.27929, 71.27931, 71.27931, 71.27928, 71.27928, 71.2793, 71.27928, 
    71.2793, 71.27927, 71.2793, 71.27927, 71.2793, 71.2793, 71.27927, 
    71.27929, 71.27927, 71.27927, 71.27929, 71.27937, 71.2794, 71.27937, 
    71.27939, 71.27939, 71.27937, 71.27937, 71.27939, 71.27938, 71.27936, 
    71.27936, 71.27938, 71.27935, 71.27937, 71.27935, 71.27937, 71.27935, 
    71.27937, 71.27934, 71.27937, 71.27937, 71.27934, 71.27937, 71.27934, 
    71.27934, 71.27936, 71.27944, 71.27946, 71.27946, 71.27944, 71.27946, 
    71.27943, 71.27943, 71.27946, 71.27946, 71.27943, 71.27945, 71.27943, 
    71.27943, 71.27945, 71.27942, 71.27944, 71.27942, 71.27944, 71.27942, 
    71.27944, 71.27943, 71.27941, 71.27943, 71.27941, 71.27943, 71.2794, 
    71.27951, 71.27953, 71.27951, 71.27953, 71.27953, 71.27951, 71.2795, 
    71.27953, 71.27953, 71.2795, 71.27953, 71.2795, 71.2795, 71.27952, 
    71.2795, 71.27952, 71.27949, 71.27951, 71.27949, 71.27951, 71.27951, 
    71.27949, 71.27951, 71.27948, 71.27948, 71.2795, 71.27959, 71.27961, 
    71.27961, 71.27958, 71.2796, 71.27958, 71.27958, 71.2796, 71.2796, 
    71.27957, 71.27957, 71.27959, 71.27957, 71.27959, 71.27959, 71.27956, 
    71.27959, 71.27956, 71.27956, 71.27959, 71.27958, 71.27956, 71.27958, 
    71.27956, 71.27958, 71.27955, 71.27966, 71.27968, 71.27968, 71.27966, 
    71.27968, 71.27965, 71.27967, 71.27965, 71.27967, 71.27965, 71.27967, 
    71.27964, 71.27966, 71.27964, 71.27964, 71.27966, 71.27963, 71.27966, 
    71.27966, 71.27963, 71.27963, 71.27966, 71.27962, 71.27965, 71.27962, 
    71.27965, 71.27973, 71.27975, 71.27975, 71.27972, 71.27975, 71.27972, 
    71.27972, 71.27975, 71.27974, 71.27972, 71.27974, 71.27972, 71.27974, 
    71.27971, 71.27973, 71.27971, 71.27973, 71.27971, 71.27972, 71.2797, 
    71.2797, 71.27972, 71.27972, 71.27969, 71.27972, 71.27969, 71.27982, 
    71.2798, 71.2798, 71.27982, 71.27982, 71.27979, 71.27982, 71.27979, 
    71.27982, 71.27979, 71.27979, 71.27981, 71.27981, 71.27979, 71.27981, 
    71.27978, 71.2798, 71.27978, 71.27978, 71.2798, 71.27977, 71.27979, 
    71.27977, 71.27979, 71.27977, 71.27979, 71.2799, 71.27987, 71.27987, 
    71.27989, 71.27987, 71.27989, 71.27988, 71.27986, 71.27986, 71.27988, 
    71.27988, 71.27985, 71.27988, 71.27985, 71.27985, 71.27988, 71.27988, 
    71.27985, 71.27987, 71.27985, 71.27985, 71.27987, 71.27984, 71.27986, 
    71.27984, 71.27985 ;

 area = 9.902211e-05, 9.902174e-05, 9.902174e-05, 9.902209e-05, 9.902172e-05, 
    9.902208e-05, 9.902207e-05, 9.902169e-05, 9.902168e-05, 9.902204e-05, 
    9.902203e-05, 9.902166e-05, 9.902201e-05, 9.902164e-05, 9.902163e-05, 
    9.902199e-05, 9.902198e-05, 9.902161e-05, 9.902196e-05, 9.902159e-05, 
    9.902158e-05, 9.902194e-05, 9.902156e-05, 9.902192e-05, 9.902155e-05, 
    4.951087e-05, 9.902174e-05, 9.902138e-05, 9.902137e-05, 9.902173e-05, 
    9.902172e-05, 9.902135e-05, 9.90217e-05, 9.902133e-05, 9.902168e-05, 
    9.902132e-05, 9.90213e-05, 9.902166e-05, 9.902164e-05, 9.902128e-05, 
    9.902163e-05, 9.902126e-05, 9.902161e-05, 9.902124e-05, 9.902123e-05, 
    9.902159e-05, 9.902121e-05, 9.902157e-05, 9.902119e-05, 9.902156e-05, 
    9.902118e-05, 9.902155e-05, 9.902102e-05, 9.902138e-05, 9.902137e-05, 
    9.9021e-05, 9.902135e-05, 9.902099e-05, 9.902097e-05, 9.902133e-05, 
    9.902132e-05, 9.902095e-05, 9.90213e-05, 9.902093e-05, 9.902128e-05, 
    9.902092e-05, 9.902126e-05, 9.90209e-05, 9.902124e-05, 9.902088e-05, 
    9.902123e-05, 9.902086e-05, 9.902084e-05, 9.902121e-05, 9.902119e-05, 
    9.902083e-05, 9.902118e-05, 9.902081e-05, 9.902065e-05, 9.902102e-05, 
    9.9021e-05, 9.902064e-05, 9.902099e-05, 9.902062e-05, 9.902097e-05, 
    9.90206e-05, 9.902095e-05, 9.902059e-05, 9.902094e-05, 9.902057e-05, 
    9.902092e-05, 9.902055e-05, 9.902054e-05, 9.90209e-05, 9.902052e-05, 
    9.902088e-05, 9.902086e-05, 9.90205e-05, 9.902048e-05, 9.902084e-05, 
    9.902046e-05, 9.902083e-05, 9.902046e-05, 9.902081e-05, 9.902029e-05, 
    9.902065e-05, 9.902064e-05, 9.902028e-05, 9.902062e-05, 9.902026e-05, 
    9.902024e-05, 9.90206e-05, 9.902059e-05, 9.902022e-05, 9.90202e-05, 
    9.902057e-05, 9.902019e-05, 9.902055e-05, 9.902054e-05, 9.902017e-05, 
    9.902052e-05, 9.902015e-05, 9.902014e-05, 9.90205e-05, 9.902048e-05, 
    9.902012e-05, 9.902046e-05, 9.90201e-05, 9.902046e-05, 9.902009e-05, 
    9.901992e-05, 9.902028e-05, 9.901991e-05, 9.902028e-05, 9.902026e-05, 
    9.901989e-05, 9.901988e-05, 9.902024e-05, 9.902022e-05, 9.901986e-05, 
    9.90202e-05, 9.901984e-05, 9.901982e-05, 9.902019e-05, 9.90198e-05, 
    9.902017e-05, 9.901979e-05, 9.902015e-05, 9.901977e-05, 9.902013e-05, 
    9.902012e-05, 9.901975e-05, 9.90201e-05, 9.901973e-05, 9.901972e-05, 
    9.902009e-05, 9.901955e-05, 9.901992e-05, 9.901991e-05, 9.901955e-05, 
    9.90199e-05, 9.901953e-05, 9.901951e-05, 9.901988e-05, 9.901986e-05, 
    9.901949e-05, 9.901984e-05, 9.901947e-05, 9.901946e-05, 9.901982e-05, 
    9.901944e-05, 9.90198e-05, 9.901942e-05, 9.901979e-05, 9.90194e-05, 
    9.901977e-05, 9.901975e-05, 9.901939e-05, 9.901974e-05, 9.901937e-05, 
    9.901972e-05, 9.901936e-05, 9.901919e-05, 9.901955e-05, 9.901918e-05, 
    9.901955e-05, 9.901953e-05, 9.901916e-05, 9.901915e-05, 9.901951e-05, 
    9.90195e-05, 9.901913e-05, 9.901911e-05, 9.901947e-05, 9.90191e-05, 
    9.901946e-05, 9.901907e-05, 9.901944e-05, 9.901906e-05, 9.901942e-05, 
    9.901904e-05, 9.90194e-05, 9.901939e-05, 9.901902e-05, 9.901937e-05, 
    9.9019e-05, 9.901899e-05, 9.901936e-05, 9.901919e-05, 9.901883e-05, 
    9.901882e-05, 9.901918e-05, 9.90188e-05, 9.901916e-05, 9.901915e-05, 
    9.901878e-05, 9.901877e-05, 9.901913e-05, 9.901911e-05, 9.901875e-05, 
    9.901873e-05, 9.90191e-05, 9.901871e-05, 9.901907e-05, 9.90187e-05, 
    9.901906e-05, 9.901867e-05, 9.901904e-05, 9.901902e-05, 9.901866e-05, 
    9.901901e-05, 9.901864e-05, 9.901863e-05, 9.901899e-05, 9.901846e-05, 
    9.901883e-05, 9.901846e-05, 9.901882e-05, 9.90188e-05, 9.901843e-05, 
    9.901842e-05, 9.901878e-05, 9.90184e-05, 9.901876e-05, 9.901838e-05, 
    9.901875e-05, 9.901873e-05, 9.901836e-05, 9.901835e-05, 9.901871e-05, 
    9.90187e-05, 9.901833e-05, 9.901867e-05, 9.901831e-05, 9.901866e-05, 
    9.90183e-05, 9.901864e-05, 9.901827e-05, 9.901863e-05, 9.901827e-05, 
    9.90181e-05, 9.901846e-05, 9.901809e-05, 9.901846e-05, 9.901843e-05, 
    9.901807e-05, 9.901842e-05, 9.901806e-05, 9.901803e-05, 9.90184e-05, 
    9.901802e-05, 9.901838e-05, 9.901837e-05, 9.9018e-05, 9.901798e-05, 
    9.901835e-05, 9.901797e-05, 9.901833e-05, 9.901795e-05, 9.901831e-05, 
    9.901793e-05, 9.90183e-05, 9.901827e-05, 9.901791e-05, 9.901827e-05, 
    9.90179e-05, 9.90181e-05, 9.901774e-05, 9.901809e-05, 9.901772e-05, 
    9.901771e-05, 9.901807e-05, 9.901769e-05, 9.901806e-05, 9.901803e-05, 
    9.901767e-05, 9.901766e-05, 9.901802e-05, 9.9018e-05, 9.901763e-05, 
    9.901798e-05, 9.901762e-05, 9.90176e-05, 9.901796e-05, 9.901758e-05, 
    9.901795e-05, 9.901757e-05, 9.901793e-05, 9.901791e-05, 9.901755e-05, 
    9.90179e-05, 9.901754e-05, 9.901774e-05, 9.901737e-05, 9.901773e-05, 
    9.901736e-05, 9.901734e-05, 9.901771e-05, 9.901733e-05, 9.901768e-05, 
    9.901731e-05, 9.901767e-05, 9.901766e-05, 9.901728e-05, 9.901727e-05, 
    9.901763e-05, 9.901762e-05, 9.901726e-05, 9.901723e-05, 9.90176e-05, 
    9.901722e-05, 9.901758e-05, 9.901757e-05, 9.90172e-05, 9.901755e-05, 
    9.901718e-05, 9.901718e-05, 9.901754e-05 ;

 topo = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0 ;

 landfrac = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 landmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 pftmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 ACTUAL_IMMOB =
  4.490659e-14, 4.502776e-14, 4.500422e-14, 4.510187e-14, 4.504772e-14, 
    4.511163e-14, 4.493118e-14, 4.503255e-14, 4.496786e-14, 4.491753e-14, 
    4.529107e-14, 4.510622e-14, 4.548291e-14, 4.536523e-14, 4.566065e-14, 
    4.546458e-14, 4.570015e-14, 4.565504e-14, 4.579087e-14, 4.575198e-14, 
    4.592545e-14, 4.580882e-14, 4.601533e-14, 4.589763e-14, 4.591603e-14, 
    4.580496e-14, 4.514348e-14, 4.526806e-14, 4.513609e-14, 4.515386e-14, 
    4.51459e-14, 4.504883e-14, 4.499986e-14, 4.489735e-14, 4.491597e-14, 
    4.499127e-14, 4.516186e-14, 4.510401e-14, 4.524983e-14, 4.524654e-14, 
    4.540864e-14, 4.533558e-14, 4.560769e-14, 4.553044e-14, 4.57536e-14, 
    4.569751e-14, 4.575096e-14, 4.573476e-14, 4.575117e-14, 4.56689e-14, 
    4.570415e-14, 4.563174e-14, 4.534926e-14, 4.543234e-14, 4.518434e-14, 
    4.503489e-14, 4.493562e-14, 4.48651e-14, 4.487507e-14, 4.489407e-14, 
    4.499171e-14, 4.508348e-14, 4.515335e-14, 4.520005e-14, 4.524606e-14, 
    4.538511e-14, 4.545872e-14, 4.562329e-14, 4.559364e-14, 4.564389e-14, 
    4.569193e-14, 4.577248e-14, 4.575923e-14, 4.57947e-14, 4.564259e-14, 
    4.57437e-14, 4.557676e-14, 4.562242e-14, 4.525843e-14, 4.511962e-14, 
    4.506046e-14, 4.500874e-14, 4.488274e-14, 4.496976e-14, 4.493546e-14, 
    4.501708e-14, 4.506889e-14, 4.504327e-14, 4.520133e-14, 4.51399e-14, 
    4.546308e-14, 4.532399e-14, 4.568633e-14, 4.559973e-14, 4.570708e-14, 
    4.565232e-14, 4.574612e-14, 4.56617e-14, 4.580791e-14, 4.583971e-14, 
    4.581798e-14, 4.590147e-14, 4.565702e-14, 4.575095e-14, 4.504255e-14, 
    4.504672e-14, 4.50662e-14, 4.498056e-14, 4.497533e-14, 4.489683e-14, 
    4.496669e-14, 4.499642e-14, 4.50719e-14, 4.51165e-14, 4.515889e-14, 
    4.525204e-14, 4.535595e-14, 4.550115e-14, 4.560534e-14, 4.567514e-14, 
    4.563236e-14, 4.567013e-14, 4.56279e-14, 4.56081e-14, 4.582779e-14, 
    4.570447e-14, 4.588947e-14, 4.587924e-14, 4.579554e-14, 4.58804e-14, 
    4.504966e-14, 4.502562e-14, 4.494205e-14, 4.500745e-14, 4.488828e-14, 
    4.495499e-14, 4.499331e-14, 4.514116e-14, 4.517365e-14, 4.520372e-14, 
    4.526313e-14, 4.533932e-14, 4.547283e-14, 4.558886e-14, 4.569473e-14, 
    4.568698e-14, 4.56897e-14, 4.571333e-14, 4.565478e-14, 4.572294e-14, 
    4.573436e-14, 4.570447e-14, 4.587787e-14, 4.582837e-14, 4.587903e-14, 
    4.58468e-14, 4.503343e-14, 4.50739e-14, 4.505203e-14, 4.509313e-14, 
    4.506417e-14, 4.519288e-14, 4.523144e-14, 4.541174e-14, 4.533781e-14, 
    4.545548e-14, 4.534978e-14, 4.536851e-14, 4.545926e-14, 4.53555e-14, 
    4.558244e-14, 4.542859e-14, 4.571425e-14, 4.556073e-14, 4.572385e-14, 
    4.569427e-14, 4.574327e-14, 4.578711e-14, 4.584228e-14, 4.594395e-14, 
    4.592042e-14, 4.600542e-14, 4.51342e-14, 4.518662e-14, 4.518203e-14, 
    4.523689e-14, 4.527743e-14, 4.536528e-14, 4.550603e-14, 4.545313e-14, 
    4.555025e-14, 4.556973e-14, 4.542219e-14, 4.551277e-14, 4.522171e-14, 
    4.526876e-14, 4.524076e-14, 4.513832e-14, 4.546528e-14, 4.529759e-14, 
    4.560706e-14, 4.551639e-14, 4.578086e-14, 4.564937e-14, 4.590746e-14, 
    4.601754e-14, 4.612116e-14, 4.624199e-14, 4.521525e-14, 4.517964e-14, 
    4.524341e-14, 4.533154e-14, 4.541332e-14, 4.552192e-14, 4.553304e-14, 
    4.555336e-14, 4.560599e-14, 4.565023e-14, 4.555976e-14, 4.566132e-14, 
    4.527962e-14, 4.547984e-14, 4.516615e-14, 4.526067e-14, 4.532636e-14, 
    4.529757e-14, 4.544709e-14, 4.548229e-14, 4.562519e-14, 4.555137e-14, 
    4.599036e-14, 4.579634e-14, 4.633398e-14, 4.618399e-14, 4.516718e-14, 
    4.521514e-14, 4.538182e-14, 4.530255e-14, 4.552917e-14, 4.558485e-14, 
    4.563014e-14, 4.568796e-14, 4.569422e-14, 4.572846e-14, 4.567234e-14, 
    4.572626e-14, 4.552215e-14, 4.56134e-14, 4.536281e-14, 4.542384e-14, 
    4.539578e-14, 4.536497e-14, 4.546003e-14, 4.556118e-14, 4.556338e-14, 
    4.559576e-14, 4.568695e-14, 4.553009e-14, 4.60153e-14, 4.571581e-14, 
    4.52674e-14, 4.53596e-14, 4.537281e-14, 4.53371e-14, 4.557929e-14, 
    4.549159e-14, 4.572763e-14, 4.566389e-14, 4.576832e-14, 4.571644e-14, 
    4.57088e-14, 4.564213e-14, 4.560059e-14, 4.549561e-14, 4.541011e-14, 
    4.534228e-14, 4.535806e-14, 4.543255e-14, 4.556737e-14, 4.569476e-14, 
    4.566686e-14, 4.576039e-14, 4.551275e-14, 4.561662e-14, 4.557649e-14, 
    4.568115e-14, 4.545171e-14, 4.5647e-14, 4.540172e-14, 4.542326e-14, 
    4.548985e-14, 4.562364e-14, 4.565328e-14, 4.568485e-14, 4.566539e-14, 
    4.55708e-14, 4.555531e-14, 4.548824e-14, 4.54697e-14, 4.541857e-14, 
    4.537621e-14, 4.54149e-14, 4.545552e-14, 4.557085e-14, 4.567464e-14, 
    4.578773e-14, 4.581541e-14, 4.594725e-14, 4.583988e-14, 4.601695e-14, 
    4.586634e-14, 4.612697e-14, 4.565836e-14, 4.586199e-14, 4.549289e-14, 
    4.553273e-14, 4.560467e-14, 4.576966e-14, 4.568066e-14, 4.578475e-14, 
    4.555471e-14, 4.54351e-14, 4.540418e-14, 4.53464e-14, 4.540551e-14, 
    4.54007e-14, 4.545723e-14, 4.543907e-14, 4.557468e-14, 4.550186e-14, 
    4.570859e-14, 4.578394e-14, 4.59965e-14, 4.612657e-14, 4.625888e-14, 
    4.631722e-14, 4.633497e-14, 4.634239e-14 ;

 AGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX_LASTYEAR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 AR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_CROP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_PEATF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BCDEP =
  8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15 ;

 BGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BTRAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BUILDHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4PROD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_DIFF_SAT =
  -1.86022e-14, -1.862564e-14, -1.862108e-14, -1.863996e-14, -1.862948e-14, 
    -1.864185e-14, -1.860694e-14, -1.862658e-14, -1.861404e-14, 
    -1.860429e-14, -1.867654e-14, -1.86408e-14, -1.871337e-14, -1.869071e-14, 
    -1.874754e-14, -1.870987e-14, -1.875512e-14, -1.874642e-14, 
    -1.877249e-14, -1.876502e-14, -1.879835e-14, -1.877593e-14, 
    -1.881552e-14, -1.879298e-14, -1.879652e-14, -1.877519e-14, 
    -1.864797e-14, -1.867211e-14, -1.864655e-14, -1.865e-14, -1.864844e-14, 
    -1.862971e-14, -1.862028e-14, -1.860038e-14, -1.860399e-14, 
    -1.861859e-14, -1.865154e-14, -1.864035e-14, -1.866847e-14, 
    -1.866783e-14, -1.869905e-14, -1.868499e-14, -1.873732e-14, 
    -1.872244e-14, -1.876534e-14, -1.875457e-14, -1.876484e-14, 
    -1.876172e-14, -1.876488e-14, -1.874909e-14, -1.875586e-14, 
    -1.874194e-14, -1.868763e-14, -1.870362e-14, -1.865587e-14, 
    -1.862707e-14, -1.860781e-14, -1.859415e-14, -1.859608e-14, 
    -1.859977e-14, -1.861867e-14, -1.863638e-14, -1.864986e-14, 
    -1.865888e-14, -1.866774e-14, -1.869461e-14, -1.870872e-14, 
    -1.874034e-14, -1.873461e-14, -1.87443e-14, -1.87535e-14, -1.876897e-14, 
    -1.876642e-14, -1.877324e-14, -1.874402e-14, -1.876346e-14, 
    -1.873135e-14, -1.874015e-14, -1.867027e-14, -1.864336e-14, -1.8632e-14, 
    -1.862196e-14, -1.859757e-14, -1.861442e-14, -1.860779e-14, 
    -1.862355e-14, -1.863357e-14, -1.862861e-14, -1.865912e-14, 
    -1.864728e-14, -1.870956e-14, -1.868278e-14, -1.875243e-14, 
    -1.873578e-14, -1.875641e-14, -1.874588e-14, -1.876392e-14, 
    -1.874769e-14, -1.877576e-14, -1.878188e-14, -1.87777e-14, -1.879369e-14, 
    -1.874679e-14, -1.876485e-14, -1.862848e-14, -1.862929e-14, 
    -1.863304e-14, -1.861652e-14, -1.86155e-14, -1.860029e-14, -1.861381e-14, 
    -1.861957e-14, -1.863414e-14, -1.864276e-14, -1.865095e-14, 
    -1.866891e-14, -1.868894e-14, -1.871685e-14, -1.873687e-14, 
    -1.875027e-14, -1.874205e-14, -1.874931e-14, -1.874119e-14, 
    -1.873738e-14, -1.87796e-14, -1.875593e-14, -1.879139e-14, -1.878943e-14, 
    -1.87734e-14, -1.878965e-14, -1.862985e-14, -1.86252e-14, -1.860905e-14, 
    -1.862169e-14, -1.859863e-14, -1.861156e-14, -1.861899e-14, 
    -1.864755e-14, -1.865378e-14, -1.86596e-14, -1.867104e-14, -1.868571e-14, 
    -1.87114e-14, -1.873371e-14, -1.875403e-14, -1.875254e-14, -1.875307e-14, 
    -1.875761e-14, -1.874637e-14, -1.875946e-14, -1.876166e-14, 
    -1.875591e-14, -1.878917e-14, -1.877968e-14, -1.878939e-14, 
    -1.878321e-14, -1.862671e-14, -1.863453e-14, -1.863031e-14, 
    -1.863826e-14, -1.863266e-14, -1.865754e-14, -1.866498e-14, 
    -1.869969e-14, -1.868543e-14, -1.870808e-14, -1.868772e-14, 
    -1.869134e-14, -1.870886e-14, -1.868882e-14, -1.87325e-14, -1.870294e-14, 
    -1.875779e-14, -1.872835e-14, -1.875963e-14, -1.875394e-14, 
    -1.876335e-14, -1.877178e-14, -1.878235e-14, -1.880185e-14, 
    -1.879733e-14, -1.88136e-14, -1.864618e-14, -1.865631e-14, -1.86554e-14, 
    -1.866598e-14, -1.86738e-14, -1.86907e-14, -1.871777e-14, -1.870759e-14, 
    -1.872625e-14, -1.873001e-14, -1.870164e-14, -1.871908e-14, 
    -1.866307e-14, -1.867217e-14, -1.866674e-14, -1.864699e-14, 
    -1.870997e-14, -1.867772e-14, -1.87372e-14, -1.871975e-14, -1.877058e-14, 
    -1.874536e-14, -1.879485e-14, -1.881598e-14, -1.883571e-14, 
    -1.885883e-14, -1.866182e-14, -1.865494e-14, -1.866723e-14, 
    -1.868425e-14, -1.869995e-14, -1.872082e-14, -1.872294e-14, 
    -1.872686e-14, -1.873698e-14, -1.874549e-14, -1.872812e-14, 
    -1.874762e-14, -1.867432e-14, -1.871275e-14, -1.865235e-14, 
    -1.867062e-14, -1.868324e-14, -1.867768e-14, -1.870642e-14, 
    -1.871319e-14, -1.87407e-14, -1.872647e-14, -1.881079e-14, -1.877359e-14, 
    -1.887632e-14, -1.884775e-14, -1.865254e-14, -1.866178e-14, 
    -1.869391e-14, -1.867864e-14, -1.87222e-14, -1.873293e-14, -1.874162e-14, 
    -1.875275e-14, -1.875394e-14, -1.876052e-14, -1.874973e-14, 
    -1.876009e-14, -1.872086e-14, -1.873841e-14, -1.869022e-14, 
    -1.870197e-14, -1.869656e-14, -1.869063e-14, -1.870891e-14, -1.87284e-14, 
    -1.872878e-14, -1.873504e-14, -1.875271e-14, -1.872237e-14, 
    -1.881564e-14, -1.875823e-14, -1.867186e-14, -1.868966e-14, 
    -1.869216e-14, -1.868527e-14, -1.873185e-14, -1.871499e-14, 
    -1.876036e-14, -1.874811e-14, -1.876816e-14, -1.875821e-14, 
    -1.875674e-14, -1.874393e-14, -1.873595e-14, -1.871577e-14, 
    -1.869934e-14, -1.868627e-14, -1.86893e-14, -1.870366e-14, -1.872958e-14, 
    -1.875406e-14, -1.874871e-14, -1.876664e-14, -1.871905e-14, 
    -1.873905e-14, -1.873133e-14, -1.875143e-14, -1.870733e-14, -1.8745e-14, 
    -1.86977e-14, -1.870185e-14, -1.871466e-14, -1.874043e-14, -1.874607e-14, 
    -1.875216e-14, -1.87484e-14, -1.873023e-14, -1.872724e-14, -1.871434e-14, 
    -1.871079e-14, -1.870094e-14, -1.86928e-14, -1.870025e-14, -1.870807e-14, 
    -1.873023e-14, -1.87502e-14, -1.87719e-14, -1.877719e-14, -1.880256e-14, 
    -1.878196e-14, -1.881597e-14, -1.878714e-14, -1.883695e-14, 
    -1.874713e-14, -1.878622e-14, -1.871523e-14, -1.872288e-14, 
    -1.873677e-14, -1.876848e-14, -1.875134e-14, -1.877136e-14, 
    -1.872712e-14, -1.870417e-14, -1.869818e-14, -1.868707e-14, 
    -1.869843e-14, -1.869751e-14, -1.870837e-14, -1.870488e-14, 
    -1.873096e-14, -1.871695e-14, -1.875672e-14, -1.87712e-14, -1.881191e-14, 
    -1.883679e-14, -1.886199e-14, -1.887311e-14, -1.887648e-14, -1.88779e-14 ;

 CH4_SURF_DIFF_UNSAT =
  1.521921e-11, 1.52148e-11, 1.521572e-11, 1.521168e-11, 1.521399e-11, 
    1.521124e-11, 1.521839e-11, 1.521461e-11, 1.521709e-11, 1.521885e-11, 
    1.520199e-11, 1.521148e-11, 1.518925e-11, 1.519746e-11, 1.508703e-11, 
    1.519061e-11, 1.508749e-11, 1.508694e-11, 1.50874e-11, 1.508764e-11, 
    1.50842e-11, 1.508719e-11, 1.507991e-11, 1.508518e-11, 1.508455e-11, 
    1.508724e-11, 1.520977e-11, 1.52033e-11, 1.521011e-11, 1.520927e-11, 
    1.520965e-11, 1.521395e-11, 1.521589e-11, 1.521952e-11, 1.52189e-11, 
    1.521622e-11, 1.520888e-11, 1.521158e-11, 1.520434e-11, 1.520452e-11, 
    1.519458e-11, 1.519933e-11, 1.508597e-11, 1.508352e-11, 1.508763e-11, 
    1.508747e-11, 1.508764e-11, 1.508764e-11, 1.508764e-11, 1.508715e-11, 
    1.508752e-11, 1.508652e-11, 1.519848e-11, 1.519294e-11, 1.520778e-11, 
    1.521451e-11, 1.521823e-11, 1.522054e-11, 1.522023e-11, 1.521962e-11, 
    1.52162e-11, 1.521249e-11, 1.52093e-11, 1.520698e-11, 1.520454e-11, 
    1.519615e-11, 1.519104e-11, 1.508633e-11, 1.50856e-11, 1.508675e-11, 
    1.508742e-11, 1.508755e-11, 1.508761e-11, 1.508736e-11, 1.508673e-11, 
    1.508764e-11, 1.508512e-11, 1.508632e-11, 1.520384e-11, 1.521088e-11, 
    1.521346e-11, 1.521555e-11, 1.521999e-11, 1.521702e-11, 1.521824e-11, 
    1.521523e-11, 1.521311e-11, 1.521418e-11, 1.520692e-11, 1.520994e-11, 
    1.519073e-11, 1.520004e-11, 1.508736e-11, 1.508577e-11, 1.508754e-11, 
    1.50869e-11, 1.508764e-11, 1.508705e-11, 1.50872e-11, 1.508667e-11, 
    1.508706e-11, 1.508505e-11, 1.508698e-11, 1.508764e-11, 1.521421e-11, 
    1.521404e-11, 1.521323e-11, 1.521662e-11, 1.521681e-11, 1.521954e-11, 
    1.521713e-11, 1.521602e-11, 1.521299e-11, 1.521102e-11, 1.520903e-11, 
    1.520421e-11, 1.519805e-11, 1.518787e-11, 1.508591e-11, 1.508723e-11, 
    1.508653e-11, 1.508717e-11, 1.508644e-11, 1.508598e-11, 1.50869e-11, 
    1.508752e-11, 1.508543e-11, 1.508573e-11, 1.508735e-11, 1.50857e-11, 
    1.521392e-11, 1.521489e-11, 1.521801e-11, 1.52156e-11, 1.521981e-11, 
    1.521755e-11, 1.521614e-11, 1.520988e-11, 1.520831e-11, 1.520679e-11, 
    1.52036e-11, 1.51991e-11, 1.519001e-11, 1.508547e-11, 1.508744e-11, 
    1.508737e-11, 1.50874e-11, 1.508757e-11, 1.508694e-11, 1.508762e-11, 
    1.508764e-11, 1.508752e-11, 1.508577e-11, 1.508689e-11, 1.508574e-11, 
    1.508653e-11, 1.521458e-11, 1.52129e-11, 1.521382e-11, 1.521206e-11, 
    1.521331e-11, 1.520734e-11, 1.520533e-11, 1.519436e-11, 1.519919e-11, 
    1.519128e-11, 1.519845e-11, 1.519725e-11, 1.5191e-11, 1.519808e-11, 
    1.508528e-11, 1.519319e-11, 1.508758e-11, 1.50846e-11, 1.508762e-11, 
    1.508744e-11, 1.508765e-11, 1.508744e-11, 1.508662e-11, 1.508347e-11, 
    1.508439e-11, 1.508047e-11, 1.52102e-11, 1.520766e-11, 1.520789e-11, 
    1.520504e-11, 1.520279e-11, 1.519746e-11, 1.51875e-11, 1.519146e-11, 
    1.508425e-11, 1.50849e-11, 1.519365e-11, 1.518697e-11, 1.520585e-11, 
    1.520328e-11, 1.520483e-11, 1.521001e-11, 1.519057e-11, 1.520162e-11, 
    1.508595e-11, 1.518669e-11, 1.508749e-11, 1.508685e-11, 1.508485e-11, 
    1.507977e-11, 1.50725e-11, 1.506074e-11, 1.520619e-11, 1.520801e-11, 
    1.520469e-11, 1.519958e-11, 1.519426e-11, 1.518625e-11, 1.508362e-11, 
    1.508436e-11, 1.508593e-11, 1.508686e-11, 1.508457e-11, 1.508704e-11, 
    1.520265e-11, 1.518949e-11, 1.520868e-11, 1.520373e-11, 1.51999e-11, 
    1.520162e-11, 1.519189e-11, 1.518931e-11, 1.508638e-11, 1.508429e-11, 
    1.508127e-11, 1.508734e-11, 1.504933e-11, 1.506683e-11, 1.520863e-11, 
    1.52062e-11, 1.519638e-11, 1.520133e-11, 1.508347e-11, 1.508535e-11, 
    1.508648e-11, 1.508738e-11, 1.508744e-11, 1.508763e-11, 1.50872e-11, 
    1.508763e-11, 1.518624e-11, 1.508611e-11, 1.519762e-11, 1.519354e-11, 
    1.519546e-11, 1.519748e-11, 1.519096e-11, 1.508462e-11, 1.508469e-11, 
    1.508566e-11, 1.508736e-11, 1.508351e-11, 1.507989e-11, 1.508758e-11, 
    1.520336e-11, 1.519782e-11, 1.519697e-11, 1.519924e-11, 1.508519e-11, 
    1.51886e-11, 1.508763e-11, 1.508708e-11, 1.508757e-11, 1.508759e-11, 
    1.508755e-11, 1.508672e-11, 1.508579e-11, 1.51883e-11, 1.519448e-11, 
    1.519892e-11, 1.519792e-11, 1.519292e-11, 1.508482e-11, 1.508744e-11, 
    1.508712e-11, 1.508761e-11, 1.518697e-11, 1.508618e-11, 1.508511e-11, 
    1.508731e-11, 1.519156e-11, 1.50868e-11, 1.519506e-11, 1.519358e-11, 
    1.518874e-11, 1.508634e-11, 1.508692e-11, 1.508735e-11, 1.50871e-11, 
    1.508493e-11, 1.508442e-11, 1.518886e-11, 1.519024e-11, 1.51939e-11, 
    1.519675e-11, 1.519415e-11, 1.519128e-11, 1.508493e-11, 1.508723e-11, 
    1.508743e-11, 1.50871e-11, 1.508331e-11, 1.508666e-11, 1.507979e-11, 
    1.508605e-11, 1.507199e-11, 1.508699e-11, 1.508617e-11, 1.518851e-11, 
    1.508361e-11, 1.508589e-11, 1.508756e-11, 1.50873e-11, 1.508745e-11, 
    1.50844e-11, 1.519274e-11, 1.519489e-11, 1.519866e-11, 1.51948e-11, 
    1.519512e-11, 1.519116e-11, 1.519247e-11, 1.508505e-11, 1.518782e-11, 
    1.508755e-11, 1.508746e-11, 1.508096e-11, 1.507204e-11, 1.505882e-11, 
    1.505158e-11, 1.50492e-11, 1.504818e-11 ;

 CH4_SURF_EBUL_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_EBUL_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_CTRUNC =
  1.931948e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 1.931948e-23, 
    1.931945e-23, 1.931947e-23, 1.931944e-23, 1.931944e-23, 1.931942e-23, 
    1.931944e-23, 1.931942e-23, 1.931942e-23, 1.931941e-23, 1.931941e-23, 
    1.93194e-23, 1.931941e-23, 1.931939e-23, 1.93194e-23, 1.93194e-23, 
    1.931941e-23, 1.931946e-23, 1.931945e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931946e-23, 1.931947e-23, 1.931945e-23, 1.931946e-23, 
    1.931944e-23, 1.931945e-23, 1.931943e-23, 1.931943e-23, 1.931941e-23, 
    1.931942e-23, 1.931941e-23, 1.931941e-23, 1.931941e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931945e-23, 1.931944e-23, 1.931946e-23, 
    1.931947e-23, 1.931948e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 
    1.931948e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 
    1.931944e-23, 1.931944e-23, 1.931942e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931941e-23, 1.931941e-23, 1.931941e-23, 1.931942e-23, 
    1.931941e-23, 1.931943e-23, 1.931942e-23, 1.931945e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 
    1.931944e-23, 1.931945e-23, 1.931942e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931941e-23, 1.931942e-23, 1.931941e-23, 1.931941e-23, 
    1.931941e-23, 1.93194e-23, 1.931942e-23, 1.931941e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931948e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 
    1.931945e-23, 1.931945e-23, 1.931943e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931943e-23, 1.931941e-23, 
    1.931942e-23, 1.93194e-23, 1.93194e-23, 1.931941e-23, 1.93194e-23, 
    1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 
    1.931948e-23, 1.931948e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 
    1.931945e-23, 1.931945e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931942e-23, 
    1.931941e-23, 1.931942e-23, 1.93194e-23, 1.931941e-23, 1.93194e-23, 
    1.931941e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931944e-23, 1.931945e-23, 
    1.931944e-23, 1.931945e-23, 1.931944e-23, 1.931944e-23, 1.931945e-23, 
    1.931943e-23, 1.931944e-23, 1.931942e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931941e-23, 1.931941e-23, 1.931941e-23, 1.93194e-23, 
    1.93194e-23, 1.931939e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931945e-23, 1.931944e-23, 1.931943e-23, 1.931944e-23, 
    1.931943e-23, 1.931943e-23, 1.931944e-23, 1.931943e-23, 1.931946e-23, 
    1.931945e-23, 1.931946e-23, 1.931946e-23, 1.931944e-23, 1.931945e-23, 
    1.931943e-23, 1.931943e-23, 1.931941e-23, 1.931942e-23, 1.93194e-23, 
    1.931939e-23, 1.931938e-23, 1.931937e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931945e-23, 1.931944e-23, 1.931943e-23, 1.931943e-23, 
    1.931943e-23, 1.931943e-23, 1.931942e-23, 1.931943e-23, 1.931942e-23, 
    1.931945e-23, 1.931944e-23, 1.931946e-23, 1.931945e-23, 1.931945e-23, 
    1.931945e-23, 1.931944e-23, 1.931944e-23, 1.931942e-23, 1.931943e-23, 
    1.931939e-23, 1.931941e-23, 1.931936e-23, 1.931938e-23, 1.931946e-23, 
    1.931946e-23, 1.931944e-23, 1.931945e-23, 1.931943e-23, 1.931943e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931941e-23, 1.931942e-23, 
    1.931941e-23, 1.931943e-23, 1.931942e-23, 1.931944e-23, 1.931944e-23, 
    1.931944e-23, 1.931944e-23, 1.931944e-23, 1.931943e-23, 1.931943e-23, 
    1.931943e-23, 1.931942e-23, 1.931943e-23, 1.931939e-23, 1.931942e-23, 
    1.931945e-23, 1.931945e-23, 1.931944e-23, 1.931945e-23, 1.931943e-23, 
    1.931944e-23, 1.931941e-23, 1.931942e-23, 1.931941e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931943e-23, 1.931944e-23, 1.931944e-23, 
    1.931945e-23, 1.931945e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931941e-23, 1.931943e-23, 1.931942e-23, 1.931943e-23, 
    1.931942e-23, 1.931944e-23, 1.931942e-23, 1.931944e-23, 1.931944e-23, 
    1.931944e-23, 1.931942e-23, 1.931942e-23, 1.931942e-23, 1.931942e-23, 
    1.931943e-23, 1.931943e-23, 1.931944e-23, 1.931944e-23, 1.931944e-23, 
    1.931944e-23, 1.931944e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931941e-23, 1.931941e-23, 1.93194e-23, 1.931941e-23, 1.931939e-23, 
    1.93194e-23, 1.931938e-23, 1.931942e-23, 1.93194e-23, 1.931944e-23, 
    1.931943e-23, 1.931943e-23, 1.931941e-23, 1.931942e-23, 1.931941e-23, 
    1.931943e-23, 1.931944e-23, 1.931944e-23, 1.931945e-23, 1.931944e-23, 
    1.931944e-23, 1.931944e-23, 1.931944e-23, 1.931943e-23, 1.931943e-23, 
    1.931942e-23, 1.931941e-23, 1.931939e-23, 1.931938e-23, 1.931937e-23, 
    1.931937e-23, 1.931936e-23, 1.931936e-23 ;

 COL_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_NTRUNC =
  1.975381e-24, 1.97538e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975381e-24, 1.97538e-24, 1.97538e-24, 1.975381e-24, 
    1.975377e-24, 1.975379e-24, 1.975374e-24, 1.975376e-24, 1.975372e-24, 
    1.975375e-24, 1.975372e-24, 1.975372e-24, 1.975371e-24, 1.975371e-24, 
    1.975369e-24, 1.975371e-24, 1.975368e-24, 1.97537e-24, 1.975369e-24, 
    1.975371e-24, 1.975378e-24, 1.975377e-24, 1.975379e-24, 1.975378e-24, 
    1.975378e-24, 1.975379e-24, 1.97538e-24, 1.975381e-24, 1.975381e-24, 
    1.97538e-24, 1.975378e-24, 1.975379e-24, 1.975377e-24, 1.975377e-24, 
    1.975375e-24, 1.975376e-24, 1.975373e-24, 1.975374e-24, 1.975371e-24, 
    1.975372e-24, 1.975371e-24, 1.975371e-24, 1.975371e-24, 1.975372e-24, 
    1.975372e-24, 1.975373e-24, 1.975376e-24, 1.975375e-24, 1.975378e-24, 
    1.97538e-24, 1.975381e-24, 1.975381e-24, 1.975381e-24, 1.975381e-24, 
    1.97538e-24, 1.975379e-24, 1.975378e-24, 1.975378e-24, 1.975377e-24, 
    1.975376e-24, 1.975375e-24, 1.975373e-24, 1.975373e-24, 1.975373e-24, 
    1.975372e-24, 1.975371e-24, 1.975371e-24, 1.975371e-24, 1.975373e-24, 
    1.975371e-24, 1.975373e-24, 1.975373e-24, 1.975377e-24, 1.975379e-24, 
    1.975379e-24, 1.97538e-24, 1.975381e-24, 1.97538e-24, 1.975381e-24, 
    1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975378e-24, 
    1.975375e-24, 1.975376e-24, 1.975372e-24, 1.975373e-24, 1.975372e-24, 
    1.975372e-24, 1.975371e-24, 1.975372e-24, 1.975371e-24, 1.97537e-24, 
    1.975371e-24, 1.97537e-24, 1.975372e-24, 1.975371e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975381e-24, 
    1.97538e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 
    1.975377e-24, 1.975376e-24, 1.975374e-24, 1.975373e-24, 1.975372e-24, 
    1.975373e-24, 1.975372e-24, 1.975373e-24, 1.975373e-24, 1.97537e-24, 
    1.975372e-24, 1.97537e-24, 1.97537e-24, 1.975371e-24, 1.97537e-24, 
    1.975379e-24, 1.97538e-24, 1.975381e-24, 1.97538e-24, 1.975381e-24, 
    1.97538e-24, 1.97538e-24, 1.975378e-24, 1.975378e-24, 1.975378e-24, 
    1.975377e-24, 1.975376e-24, 1.975375e-24, 1.975373e-24, 1.975372e-24, 
    1.975372e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 
    1.975371e-24, 1.975372e-24, 1.97537e-24, 1.97537e-24, 1.97537e-24, 
    1.97537e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975378e-24, 1.975377e-24, 1.975375e-24, 1.975376e-24, 
    1.975375e-24, 1.975376e-24, 1.975376e-24, 1.975375e-24, 1.975376e-24, 
    1.975373e-24, 1.975375e-24, 1.975372e-24, 1.975374e-24, 1.975372e-24, 
    1.975372e-24, 1.975371e-24, 1.975371e-24, 1.97537e-24, 1.975369e-24, 
    1.975369e-24, 1.975368e-24, 1.975379e-24, 1.975378e-24, 1.975378e-24, 
    1.975377e-24, 1.975377e-24, 1.975376e-24, 1.975374e-24, 1.975375e-24, 
    1.975374e-24, 1.975373e-24, 1.975375e-24, 1.975374e-24, 1.975378e-24, 
    1.975377e-24, 1.975377e-24, 1.975378e-24, 1.975375e-24, 1.975377e-24, 
    1.975373e-24, 1.975374e-24, 1.975371e-24, 1.975372e-24, 1.975369e-24, 
    1.975368e-24, 1.975367e-24, 1.975365e-24, 1.975378e-24, 1.975378e-24, 
    1.975377e-24, 1.975376e-24, 1.975375e-24, 1.975374e-24, 1.975374e-24, 
    1.975374e-24, 1.975373e-24, 1.975372e-24, 1.975374e-24, 1.975372e-24, 
    1.975377e-24, 1.975374e-24, 1.975378e-24, 1.975377e-24, 1.975376e-24, 
    1.975377e-24, 1.975375e-24, 1.975374e-24, 1.975373e-24, 1.975374e-24, 
    1.975368e-24, 1.975371e-24, 1.975365e-24, 1.975366e-24, 1.975378e-24, 
    1.975378e-24, 1.975376e-24, 1.975377e-24, 1.975374e-24, 1.975373e-24, 
    1.975373e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 
    1.975372e-24, 1.975374e-24, 1.975373e-24, 1.975376e-24, 1.975375e-24, 
    1.975375e-24, 1.975376e-24, 1.975375e-24, 1.975374e-24, 1.975374e-24, 
    1.975373e-24, 1.975372e-24, 1.975374e-24, 1.975368e-24, 1.975372e-24, 
    1.975377e-24, 1.975376e-24, 1.975376e-24, 1.975376e-24, 1.975373e-24, 
    1.975374e-24, 1.975372e-24, 1.975372e-24, 1.975371e-24, 1.975372e-24, 
    1.975372e-24, 1.975373e-24, 1.975373e-24, 1.975374e-24, 1.975375e-24, 
    1.975376e-24, 1.975376e-24, 1.975375e-24, 1.975373e-24, 1.975372e-24, 
    1.975372e-24, 1.975371e-24, 1.975374e-24, 1.975373e-24, 1.975373e-24, 
    1.975372e-24, 1.975375e-24, 1.975373e-24, 1.975375e-24, 1.975375e-24, 
    1.975374e-24, 1.975373e-24, 1.975372e-24, 1.975372e-24, 1.975372e-24, 
    1.975373e-24, 1.975374e-24, 1.975374e-24, 1.975375e-24, 1.975375e-24, 
    1.975376e-24, 1.975375e-24, 1.975375e-24, 1.975373e-24, 1.975372e-24, 
    1.975371e-24, 1.975371e-24, 1.975369e-24, 1.97537e-24, 1.975368e-24, 
    1.97537e-24, 1.975367e-24, 1.975372e-24, 1.97537e-24, 1.975374e-24, 
    1.975374e-24, 1.975373e-24, 1.975371e-24, 1.975372e-24, 1.975371e-24, 
    1.975374e-24, 1.975375e-24, 1.975375e-24, 1.975376e-24, 1.975375e-24, 
    1.975375e-24, 1.975375e-24, 1.975375e-24, 1.975373e-24, 1.975374e-24, 
    1.975372e-24, 1.975371e-24, 1.975368e-24, 1.975367e-24, 1.975365e-24, 
    1.975365e-24, 1.975365e-24, 1.975364e-24 ;

 CONC_CH4_SAT =
  8.381706e-08, 8.392507e-08, 8.390406e-08, 8.399109e-08, 8.394279e-08, 
    8.399978e-08, 8.383892e-08, 8.392941e-08, 8.387163e-08, 8.382672e-08, 
    8.415965e-08, 8.399495e-08, 8.432947e-08, 8.422502e-08, 8.4487e-08, 
    8.431331e-08, 8.452193e-08, 8.448185e-08, 8.460201e-08, 8.456762e-08, 
    8.472121e-08, 8.461788e-08, 8.480038e-08, 8.469648e-08, 8.471281e-08, 
    8.461448e-08, 8.402802e-08, 8.413923e-08, 8.402145e-08, 8.403732e-08, 
    8.403018e-08, 8.394383e-08, 8.390034e-08, 8.380871e-08, 8.382533e-08, 
    8.389258e-08, 8.404446e-08, 8.399287e-08, 8.41225e-08, 8.411957e-08, 
    8.426349e-08, 8.419866e-08, 8.443991e-08, 8.437134e-08, 8.456905e-08, 
    8.451944e-08, 8.456675e-08, 8.455239e-08, 8.456693e-08, 8.449414e-08, 
    8.452535e-08, 8.44612e-08, 8.421083e-08, 8.428455e-08, 8.406439e-08, 
    8.393165e-08, 8.384292e-08, 8.377995e-08, 8.378886e-08, 8.380587e-08, 
    8.389297e-08, 8.397461e-08, 8.403674e-08, 8.407828e-08, 8.411915e-08, 
    8.424295e-08, 8.430804e-08, 8.445382e-08, 8.442741e-08, 8.447206e-08, 
    8.45145e-08, 8.458581e-08, 8.457406e-08, 8.460547e-08, 8.44708e-08, 
    8.45604e-08, 8.441239e-08, 8.445294e-08, 8.413072e-08, 8.400677e-08, 
    8.395438e-08, 8.390812e-08, 8.379572e-08, 8.38734e-08, 8.38428e-08, 
    8.391545e-08, 8.396162e-08, 8.393877e-08, 8.407942e-08, 8.402481e-08, 
    8.43119e-08, 8.418847e-08, 8.450955e-08, 8.443283e-08, 8.45279e-08, 
    8.447939e-08, 8.456251e-08, 8.448771e-08, 8.461712e-08, 8.46453e-08, 
    8.462606e-08, 8.469977e-08, 8.448357e-08, 8.456679e-08, 8.393815e-08, 
    8.394188e-08, 8.395921e-08, 8.388303e-08, 8.387834e-08, 8.380827e-08, 
    8.387058e-08, 8.389713e-08, 8.396426e-08, 8.4004e-08, 8.404172e-08, 
    8.412452e-08, 8.421686e-08, 8.434553e-08, 8.443781e-08, 8.44996e-08, 
    8.44617e-08, 8.449517e-08, 8.445777e-08, 8.44402e-08, 8.463478e-08, 
    8.452567e-08, 8.468918e-08, 8.468013e-08, 8.460623e-08, 8.468115e-08, 
    8.39445e-08, 8.392305e-08, 8.384863e-08, 8.390688e-08, 8.380063e-08, 
    8.386019e-08, 8.389443e-08, 8.402606e-08, 8.40548e-08, 8.408159e-08, 
    8.413434e-08, 8.420199e-08, 8.432043e-08, 8.442326e-08, 8.451695e-08, 
    8.451008e-08, 8.45125e-08, 8.453345e-08, 8.44816e-08, 8.454195e-08, 
    8.455211e-08, 8.45256e-08, 8.467892e-08, 8.463518e-08, 8.467994e-08, 
    8.465145e-08, 8.393e-08, 8.396607e-08, 8.39466e-08, 8.398324e-08, 
    8.395746e-08, 8.407208e-08, 8.410638e-08, 8.426639e-08, 8.420068e-08, 
    8.430509e-08, 8.421126e-08, 8.422792e-08, 8.430868e-08, 8.42163e-08, 
    8.441769e-08, 8.42814e-08, 8.453426e-08, 8.439854e-08, 8.454276e-08, 
    8.451654e-08, 8.45599e-08, 8.459875e-08, 8.464748e-08, 8.473738e-08, 
    8.471656e-08, 8.479155e-08, 8.401973e-08, 8.406644e-08, 8.406225e-08, 
    8.411102e-08, 8.414708e-08, 8.422499e-08, 8.434978e-08, 8.430287e-08, 
    8.43889e-08, 8.440621e-08, 8.427542e-08, 8.43558e-08, 8.409761e-08, 
    8.413953e-08, 8.411452e-08, 8.402347e-08, 8.43138e-08, 8.416511e-08, 
    8.443935e-08, 8.435892e-08, 8.459322e-08, 8.447695e-08, 8.470511e-08, 
    8.480249e-08, 8.489351e-08, 8.500008e-08, 8.409182e-08, 8.406012e-08, 
    8.411679e-08, 8.419523e-08, 8.426763e-08, 8.436385e-08, 8.437364e-08, 
    8.43917e-08, 8.443833e-08, 8.447755e-08, 8.439749e-08, 8.448737e-08, 
    8.414941e-08, 8.432664e-08, 8.40482e-08, 8.413237e-08, 8.419057e-08, 
    8.416496e-08, 8.429748e-08, 8.432869e-08, 8.445548e-08, 8.438989e-08, 
    8.477856e-08, 8.460707e-08, 8.508074e-08, 8.4949e-08, 8.404906e-08, 
    8.409167e-08, 8.423977e-08, 8.416936e-08, 8.437021e-08, 8.441966e-08, 
    8.445973e-08, 8.451104e-08, 8.451651e-08, 8.454687e-08, 8.449712e-08, 
    8.454487e-08, 8.436405e-08, 8.444493e-08, 8.422277e-08, 8.427696e-08, 
    8.425201e-08, 8.422469e-08, 8.430897e-08, 8.439878e-08, 8.440055e-08, 
    8.442937e-08, 8.451074e-08, 8.437102e-08, 8.48009e-08, 8.45362e-08, 
    8.41381e-08, 8.422016e-08, 8.423169e-08, 8.419997e-08, 8.441471e-08, 
    8.433698e-08, 8.454611e-08, 8.448964e-08, 8.458208e-08, 8.453619e-08, 
    8.452944e-08, 8.447037e-08, 8.443359e-08, 8.434057e-08, 8.42648e-08, 
    8.420455e-08, 8.421856e-08, 8.428471e-08, 8.440423e-08, 8.451707e-08, 
    8.44924e-08, 8.457506e-08, 8.435568e-08, 8.444788e-08, 8.44123e-08, 
    8.450496e-08, 8.430165e-08, 8.447525e-08, 8.425727e-08, 8.427638e-08, 
    8.433543e-08, 8.445421e-08, 8.448026e-08, 8.450829e-08, 8.449096e-08, 
    8.440725e-08, 8.439345e-08, 8.433397e-08, 8.431761e-08, 8.427221e-08, 
    8.423465e-08, 8.4269e-08, 8.430508e-08, 8.440723e-08, 8.449926e-08, 
    8.459932e-08, 8.462371e-08, 8.47406e-08, 8.464567e-08, 8.480239e-08, 
    8.466947e-08, 8.489913e-08, 8.448509e-08, 8.466528e-08, 8.433808e-08, 
    8.437335e-08, 8.443737e-08, 8.45835e-08, 8.450453e-08, 8.459681e-08, 
    8.43929e-08, 8.428706e-08, 8.425947e-08, 8.420825e-08, 8.426064e-08, 
    8.425638e-08, 8.430647e-08, 8.429038e-08, 8.441062e-08, 8.434602e-08, 
    8.45293e-08, 8.459605e-08, 8.478375e-08, 8.489847e-08, 8.501468e-08, 
    8.506595e-08, 8.508152e-08, 8.508805e-08,
  2.311746e-10, 2.317738e-10, 2.316571e-10, 2.321405e-10, 2.318721e-10, 
    2.321888e-10, 2.312957e-10, 2.317979e-10, 2.314772e-10, 2.31228e-10, 
    2.330786e-10, 2.32162e-10, 2.340256e-10, 2.334427e-10, 2.349058e-10, 
    2.339355e-10, 2.351012e-10, 2.34877e-10, 2.355495e-10, 2.353568e-10, 
    2.362179e-10, 2.356383e-10, 2.366622e-10, 2.36079e-10, 2.361707e-10, 
    2.356193e-10, 2.323457e-10, 2.329649e-10, 2.323092e-10, 2.323975e-10, 
    2.323577e-10, 2.31878e-10, 2.316366e-10, 2.311282e-10, 2.312204e-10, 
    2.315934e-10, 2.324372e-10, 2.321503e-10, 2.328713e-10, 2.32855e-10, 
    2.336572e-10, 2.332957e-10, 2.346424e-10, 2.342594e-10, 2.353649e-10, 
    2.350872e-10, 2.35352e-10, 2.352716e-10, 2.35353e-10, 2.349457e-10, 
    2.351203e-10, 2.347614e-10, 2.333636e-10, 2.337748e-10, 2.325481e-10, 
    2.318105e-10, 2.313179e-10, 2.309688e-10, 2.310182e-10, 2.311125e-10, 
    2.315956e-10, 2.320488e-10, 2.323942e-10, 2.326253e-10, 2.328527e-10, 
    2.335429e-10, 2.33906e-10, 2.347203e-10, 2.345726e-10, 2.348222e-10, 
    2.350595e-10, 2.354587e-10, 2.353929e-10, 2.355689e-10, 2.348151e-10, 
    2.353165e-10, 2.344886e-10, 2.347153e-10, 2.329175e-10, 2.322276e-10, 
    2.319367e-10, 2.316797e-10, 2.310562e-10, 2.31487e-10, 2.313173e-10, 
    2.317203e-10, 2.319767e-10, 2.318498e-10, 2.326316e-10, 2.323279e-10, 
    2.339275e-10, 2.33239e-10, 2.350319e-10, 2.346028e-10, 2.351345e-10, 
    2.348631e-10, 2.353283e-10, 2.349097e-10, 2.356341e-10, 2.357921e-10, 
    2.356842e-10, 2.360974e-10, 2.348865e-10, 2.353523e-10, 2.318464e-10, 
    2.318671e-10, 2.319633e-10, 2.315405e-10, 2.315144e-10, 2.311258e-10, 
    2.314714e-10, 2.316187e-10, 2.319913e-10, 2.322122e-10, 2.324219e-10, 
    2.328826e-10, 2.333972e-10, 2.341153e-10, 2.346307e-10, 2.349762e-10, 
    2.347642e-10, 2.349514e-10, 2.347422e-10, 2.34644e-10, 2.357331e-10, 
    2.351221e-10, 2.36038e-10, 2.359873e-10, 2.355732e-10, 2.35993e-10, 
    2.318816e-10, 2.317625e-10, 2.313496e-10, 2.316727e-10, 2.310834e-10, 
    2.314137e-10, 2.316038e-10, 2.323349e-10, 2.324947e-10, 2.326437e-10, 
    2.329373e-10, 2.333142e-10, 2.33975e-10, 2.345494e-10, 2.350732e-10, 
    2.350348e-10, 2.350483e-10, 2.351656e-10, 2.348755e-10, 2.352132e-10, 
    2.352701e-10, 2.351217e-10, 2.359805e-10, 2.357353e-10, 2.359862e-10, 
    2.358265e-10, 2.318011e-10, 2.320014e-10, 2.318932e-10, 2.320968e-10, 
    2.319536e-10, 2.325909e-10, 2.327818e-10, 2.336735e-10, 2.33307e-10, 
    2.338894e-10, 2.333659e-10, 2.334589e-10, 2.339096e-10, 2.33394e-10, 
    2.345183e-10, 2.337573e-10, 2.351702e-10, 2.344115e-10, 2.352177e-10, 
    2.350709e-10, 2.353136e-10, 2.355312e-10, 2.358042e-10, 2.363085e-10, 
    2.361916e-10, 2.366126e-10, 2.322996e-10, 2.325595e-10, 2.325361e-10, 
    2.328075e-10, 2.330082e-10, 2.334425e-10, 2.341389e-10, 2.338769e-10, 
    2.343574e-10, 2.344541e-10, 2.337238e-10, 2.341726e-10, 2.327329e-10, 
    2.329663e-10, 2.328269e-10, 2.323205e-10, 2.339381e-10, 2.331088e-10, 
    2.346393e-10, 2.3419e-10, 2.355003e-10, 2.348496e-10, 2.361275e-10, 
    2.366742e-10, 2.371855e-10, 2.377854e-10, 2.327006e-10, 2.325242e-10, 
    2.328396e-10, 2.332766e-10, 2.336803e-10, 2.342175e-10, 2.342722e-10, 
    2.34373e-10, 2.346336e-10, 2.348529e-10, 2.344055e-10, 2.349077e-10, 
    2.330215e-10, 2.340098e-10, 2.32458e-10, 2.329265e-10, 2.332506e-10, 
    2.331079e-10, 2.338469e-10, 2.340211e-10, 2.347295e-10, 2.343629e-10, 
    2.365398e-10, 2.355779e-10, 2.382398e-10, 2.374978e-10, 2.324627e-10, 
    2.326998e-10, 2.335249e-10, 2.331324e-10, 2.342531e-10, 2.345293e-10, 
    2.347532e-10, 2.350402e-10, 2.350708e-10, 2.352407e-10, 2.349623e-10, 
    2.352295e-10, 2.342186e-10, 2.346705e-10, 2.3343e-10, 2.337324e-10, 
    2.335931e-10, 2.334407e-10, 2.339109e-10, 2.344127e-10, 2.344225e-10, 
    2.345836e-10, 2.350389e-10, 2.342576e-10, 2.366655e-10, 2.351813e-10, 
    2.329582e-10, 2.334156e-10, 2.334799e-10, 2.333029e-10, 2.345016e-10, 
    2.340674e-10, 2.352364e-10, 2.349205e-10, 2.354378e-10, 2.351809e-10, 
    2.351431e-10, 2.348127e-10, 2.346071e-10, 2.340875e-10, 2.336645e-10, 
    2.333285e-10, 2.334066e-10, 2.337756e-10, 2.344432e-10, 2.35074e-10, 
    2.34936e-10, 2.353985e-10, 2.341719e-10, 2.34687e-10, 2.344882e-10, 
    2.350062e-10, 2.338702e-10, 2.348404e-10, 2.336225e-10, 2.337291e-10, 
    2.340588e-10, 2.347225e-10, 2.34868e-10, 2.350249e-10, 2.349279e-10, 
    2.3446e-10, 2.343829e-10, 2.340506e-10, 2.339593e-10, 2.337058e-10, 
    2.334963e-10, 2.33688e-10, 2.338894e-10, 2.344598e-10, 2.349743e-10, 
    2.355345e-10, 2.35671e-10, 2.363267e-10, 2.357943e-10, 2.366739e-10, 
    2.35928e-10, 2.372174e-10, 2.348952e-10, 2.359043e-10, 2.340735e-10, 
    2.342706e-10, 2.346283e-10, 2.35446e-10, 2.350037e-10, 2.355204e-10, 
    2.343798e-10, 2.337888e-10, 2.336348e-10, 2.333491e-10, 2.336413e-10, 
    2.336175e-10, 2.33897e-10, 2.338072e-10, 2.344787e-10, 2.341179e-10, 
    2.351424e-10, 2.355161e-10, 2.365688e-10, 2.372135e-10, 2.378675e-10, 
    2.381564e-10, 2.382441e-10, 2.382809e-10,
  1.303421e-13, 1.307934e-13, 1.307055e-13, 1.310699e-13, 1.308676e-13, 
    1.311063e-13, 1.304333e-13, 1.308116e-13, 1.305699e-13, 1.303823e-13, 
    1.317779e-13, 1.310861e-13, 1.32505e-13, 1.320529e-13, 1.331893e-13, 
    1.324349e-13, 1.333413e-13, 1.331668e-13, 1.336902e-13, 1.335402e-13, 
    1.342109e-13, 1.337594e-13, 1.345574e-13, 1.341027e-13, 1.341741e-13, 
    1.337446e-13, 1.312247e-13, 1.31692e-13, 1.311972e-13, 1.312638e-13, 
    1.312338e-13, 1.30872e-13, 1.306901e-13, 1.303071e-13, 1.303765e-13, 
    1.306575e-13, 1.312937e-13, 1.310773e-13, 1.316214e-13, 1.316091e-13, 
    1.322188e-13, 1.319418e-13, 1.329845e-13, 1.326867e-13, 1.335465e-13, 
    1.333304e-13, 1.335364e-13, 1.334738e-13, 1.335372e-13, 1.332203e-13, 
    1.333561e-13, 1.33077e-13, 1.319931e-13, 1.323101e-13, 1.313773e-13, 
    1.308211e-13, 1.3045e-13, 1.301871e-13, 1.302243e-13, 1.302953e-13, 
    1.306592e-13, 1.310008e-13, 1.312613e-13, 1.314356e-13, 1.316073e-13, 
    1.321299e-13, 1.32412e-13, 1.33045e-13, 1.329302e-13, 1.331242e-13, 
    1.333088e-13, 1.336195e-13, 1.335683e-13, 1.337053e-13, 1.331187e-13, 
    1.335088e-13, 1.328649e-13, 1.330411e-13, 1.316562e-13, 1.311356e-13, 
    1.309162e-13, 1.307225e-13, 1.302529e-13, 1.305774e-13, 1.304495e-13, 
    1.307532e-13, 1.309464e-13, 1.308507e-13, 1.314404e-13, 1.312112e-13, 
    1.324287e-13, 1.31899e-13, 1.332873e-13, 1.329537e-13, 1.333672e-13, 
    1.331561e-13, 1.33518e-13, 1.331923e-13, 1.337561e-13, 1.338791e-13, 
    1.337951e-13, 1.34117e-13, 1.331743e-13, 1.335366e-13, 1.308482e-13, 
    1.308638e-13, 1.309363e-13, 1.306176e-13, 1.30598e-13, 1.303053e-13, 
    1.305656e-13, 1.306766e-13, 1.309574e-13, 1.31124e-13, 1.312822e-13, 
    1.316299e-13, 1.320185e-13, 1.325747e-13, 1.329753e-13, 1.33244e-13, 
    1.330791e-13, 1.332247e-13, 1.33062e-13, 1.329857e-13, 1.338332e-13, 
    1.333575e-13, 1.340707e-13, 1.340312e-13, 1.337086e-13, 1.340356e-13, 
    1.308747e-13, 1.307849e-13, 1.304738e-13, 1.307173e-13, 1.302734e-13, 
    1.305222e-13, 1.306653e-13, 1.312165e-13, 1.313371e-13, 1.314496e-13, 
    1.316712e-13, 1.319558e-13, 1.324657e-13, 1.329122e-13, 1.333195e-13, 
    1.332896e-13, 1.333001e-13, 1.333914e-13, 1.331657e-13, 1.334284e-13, 
    1.334727e-13, 1.333572e-13, 1.340259e-13, 1.338349e-13, 1.340304e-13, 
    1.339059e-13, 1.30814e-13, 1.30965e-13, 1.308835e-13, 1.31037e-13, 
    1.30929e-13, 1.314097e-13, 1.315538e-13, 1.322314e-13, 1.319503e-13, 
    1.323992e-13, 1.319949e-13, 1.320651e-13, 1.324149e-13, 1.320161e-13, 
    1.32888e-13, 1.322965e-13, 1.333949e-13, 1.328049e-13, 1.334319e-13, 
    1.333177e-13, 1.335066e-13, 1.336759e-13, 1.338886e-13, 1.342816e-13, 
    1.341905e-13, 1.345187e-13, 1.311899e-13, 1.31386e-13, 1.313683e-13, 
    1.315732e-13, 1.317247e-13, 1.320527e-13, 1.325931e-13, 1.323895e-13, 
    1.327629e-13, 1.328381e-13, 1.322705e-13, 1.326193e-13, 1.315168e-13, 
    1.316931e-13, 1.315878e-13, 1.312056e-13, 1.32437e-13, 1.318007e-13, 
    1.32982e-13, 1.326328e-13, 1.336519e-13, 1.331455e-13, 1.341404e-13, 
    1.345667e-13, 1.349659e-13, 1.354345e-13, 1.314925e-13, 1.313594e-13, 
    1.315974e-13, 1.319275e-13, 1.322367e-13, 1.326542e-13, 1.326967e-13, 
    1.327751e-13, 1.329776e-13, 1.331481e-13, 1.328003e-13, 1.331908e-13, 
    1.317348e-13, 1.324927e-13, 1.313094e-13, 1.31663e-13, 1.319078e-13, 
    1.318e-13, 1.323661e-13, 1.325015e-13, 1.330522e-13, 1.327672e-13, 
    1.344619e-13, 1.337123e-13, 1.357898e-13, 1.352098e-13, 1.313129e-13, 
    1.314918e-13, 1.32116e-13, 1.318185e-13, 1.326818e-13, 1.328965e-13, 
    1.330706e-13, 1.332938e-13, 1.333176e-13, 1.334498e-13, 1.332332e-13, 
    1.334411e-13, 1.326551e-13, 1.330063e-13, 1.320433e-13, 1.322772e-13, 
    1.32169e-13, 1.320514e-13, 1.324159e-13, 1.328059e-13, 1.328135e-13, 
    1.329387e-13, 1.332928e-13, 1.326854e-13, 1.345599e-13, 1.334036e-13, 
    1.31687e-13, 1.320325e-13, 1.32081e-13, 1.319473e-13, 1.32875e-13, 
    1.325375e-13, 1.334465e-13, 1.332007e-13, 1.336033e-13, 1.334033e-13, 
    1.333739e-13, 1.331169e-13, 1.32957e-13, 1.325531e-13, 1.322245e-13, 
    1.319666e-13, 1.320256e-13, 1.323108e-13, 1.328296e-13, 1.333201e-13, 
    1.332127e-13, 1.335727e-13, 1.326187e-13, 1.330191e-13, 1.328646e-13, 
    1.332673e-13, 1.323842e-13, 1.331383e-13, 1.321918e-13, 1.322746e-13, 
    1.325308e-13, 1.330467e-13, 1.331598e-13, 1.332819e-13, 1.332064e-13, 
    1.328426e-13, 1.327827e-13, 1.325244e-13, 1.324535e-13, 1.322565e-13, 
    1.320938e-13, 1.322426e-13, 1.323991e-13, 1.328425e-13, 1.332426e-13, 
    1.336785e-13, 1.337848e-13, 1.342958e-13, 1.338808e-13, 1.345665e-13, 
    1.33985e-13, 1.349908e-13, 1.33181e-13, 1.339665e-13, 1.325423e-13, 
    1.326954e-13, 1.329735e-13, 1.336096e-13, 1.332654e-13, 1.336675e-13, 
    1.327803e-13, 1.32321e-13, 1.322013e-13, 1.319822e-13, 1.322064e-13, 
    1.321879e-13, 1.324051e-13, 1.323353e-13, 1.328572e-13, 1.325768e-13, 
    1.333733e-13, 1.336642e-13, 1.344845e-13, 1.349877e-13, 1.354987e-13, 
    1.357246e-13, 1.357933e-13, 1.35822e-13,
  1.914839e-17, 1.922371e-17, 1.920904e-17, 1.926988e-17, 1.923609e-17, 
    1.927596e-17, 1.916361e-17, 1.922674e-17, 1.918641e-17, 1.915511e-17, 
    1.938865e-17, 1.927258e-17, 1.951496e-17, 1.943641e-17, 1.963394e-17, 
    1.950277e-17, 1.966039e-17, 1.963004e-17, 1.972115e-17, 1.969503e-17, 
    1.981188e-17, 1.97332e-17, 1.987232e-17, 1.979303e-17, 1.980547e-17, 
    1.973063e-17, 1.929574e-17, 1.937381e-17, 1.929114e-17, 1.930226e-17, 
    1.929725e-17, 1.923682e-17, 1.920645e-17, 1.914257e-17, 1.915415e-17, 
    1.920103e-17, 1.930726e-17, 1.927112e-17, 1.936203e-17, 1.935998e-17, 
    1.946522e-17, 1.941714e-17, 1.959832e-17, 1.954656e-17, 1.969612e-17, 
    1.96585e-17, 1.969437e-17, 1.968348e-17, 1.969452e-17, 1.963934e-17, 
    1.966298e-17, 1.961441e-17, 1.942604e-17, 1.948109e-17, 1.932124e-17, 
    1.922831e-17, 1.91664e-17, 1.912256e-17, 1.912876e-17, 1.914059e-17, 
    1.92013e-17, 1.925833e-17, 1.930185e-17, 1.933098e-17, 1.935968e-17, 
    1.944977e-17, 1.949879e-17, 1.960884e-17, 1.958888e-17, 1.962263e-17, 
    1.965476e-17, 1.970884e-17, 1.969992e-17, 1.972378e-17, 1.962168e-17, 
    1.968955e-17, 1.957753e-17, 1.960817e-17, 1.936782e-17, 1.928085e-17, 
    1.92442e-17, 1.921187e-17, 1.913353e-17, 1.918764e-17, 1.916631e-17, 
    1.921699e-17, 1.924926e-17, 1.923328e-17, 1.933178e-17, 1.929349e-17, 
    1.95017e-17, 1.940969e-17, 1.965101e-17, 1.959297e-17, 1.966491e-17, 
    1.962818e-17, 1.969116e-17, 1.963447e-17, 1.973263e-17, 1.975406e-17, 
    1.973942e-17, 1.979553e-17, 1.963134e-17, 1.969441e-17, 1.923285e-17, 
    1.923546e-17, 1.924756e-17, 1.919437e-17, 1.919109e-17, 1.914227e-17, 
    1.918568e-17, 1.92042e-17, 1.92511e-17, 1.927891e-17, 1.930534e-17, 
    1.936346e-17, 1.943044e-17, 1.952708e-17, 1.959674e-17, 1.964348e-17, 
    1.961479e-17, 1.964012e-17, 1.961182e-17, 1.959854e-17, 1.974605e-17, 
    1.966322e-17, 1.978746e-17, 1.978057e-17, 1.972436e-17, 1.978134e-17, 
    1.923728e-17, 1.922229e-17, 1.917038e-17, 1.9211e-17, 1.913695e-17, 
    1.917844e-17, 1.920232e-17, 1.929436e-17, 1.931451e-17, 1.933331e-17, 
    1.937036e-17, 1.941957e-17, 1.950813e-17, 1.958575e-17, 1.965661e-17, 
    1.965141e-17, 1.965325e-17, 1.966912e-17, 1.962985e-17, 1.967557e-17, 
    1.968327e-17, 1.966317e-17, 1.977965e-17, 1.974635e-17, 1.978042e-17, 
    1.975873e-17, 1.922716e-17, 1.925237e-17, 1.923875e-17, 1.926438e-17, 
    1.924635e-17, 1.932663e-17, 1.935072e-17, 1.946741e-17, 1.941861e-17, 
    1.949656e-17, 1.942635e-17, 1.943853e-17, 1.949927e-17, 1.943003e-17, 
    1.958153e-17, 1.947871e-17, 1.966974e-17, 1.956708e-17, 1.967618e-17, 
    1.965631e-17, 1.968918e-17, 1.971867e-17, 1.975572e-17, 1.982421e-17, 
    1.980833e-17, 1.986558e-17, 1.928993e-17, 1.932268e-17, 1.931973e-17, 
    1.935397e-17, 1.937946e-17, 1.943639e-17, 1.953028e-17, 1.949489e-17, 
    1.95598e-17, 1.957287e-17, 1.947421e-17, 1.953483e-17, 1.934455e-17, 
    1.937401e-17, 1.935643e-17, 1.929255e-17, 1.950314e-17, 1.939263e-17, 
    1.95979e-17, 1.953719e-17, 1.971447e-17, 1.962633e-17, 1.97996e-17, 
    1.987394e-17, 1.994363e-17, 2.00255e-17, 1.934049e-17, 1.931824e-17, 
    1.935802e-17, 1.941463e-17, 1.946834e-17, 1.95409e-17, 1.954829e-17, 
    1.956192e-17, 1.959713e-17, 1.962679e-17, 1.956629e-17, 1.963421e-17, 
    1.938117e-17, 1.951282e-17, 1.930988e-17, 1.936898e-17, 1.941123e-17, 
    1.939252e-17, 1.949083e-17, 1.951436e-17, 1.961009e-17, 1.956055e-17, 
    1.985565e-17, 1.972499e-17, 2.008765e-17, 1.998623e-17, 1.931048e-17, 
    1.934038e-17, 1.944737e-17, 1.939573e-17, 1.954571e-17, 1.958302e-17, 
    1.961331e-17, 1.965214e-17, 1.965628e-17, 1.967929e-17, 1.96416e-17, 
    1.967778e-17, 1.954106e-17, 1.960212e-17, 1.943476e-17, 1.947537e-17, 
    1.945658e-17, 1.943616e-17, 1.949948e-17, 1.956726e-17, 1.95686e-17, 
    1.959036e-17, 1.965191e-17, 1.954632e-17, 1.987272e-17, 1.96712e-17, 
    1.937301e-17, 1.943286e-17, 1.94413e-17, 1.941809e-17, 1.957928e-17, 
    1.952062e-17, 1.967872e-17, 1.963594e-17, 1.970601e-17, 1.96712e-17, 
    1.966608e-17, 1.962135e-17, 1.959355e-17, 1.952333e-17, 1.946621e-17, 
    1.942144e-17, 1.943168e-17, 1.948121e-17, 1.957138e-17, 1.965671e-17, 
    1.963802e-17, 1.970068e-17, 1.953474e-17, 1.960434e-17, 1.957747e-17, 
    1.964754e-17, 1.949397e-17, 1.962505e-17, 1.946054e-17, 1.947493e-17, 
    1.951945e-17, 1.960914e-17, 1.962883e-17, 1.965006e-17, 1.963694e-17, 
    1.957365e-17, 1.956324e-17, 1.951834e-17, 1.950601e-17, 1.947179e-17, 
    1.944352e-17, 1.946937e-17, 1.949656e-17, 1.957363e-17, 1.964322e-17, 
    1.971911e-17, 1.973764e-17, 1.982666e-17, 1.975434e-17, 1.987386e-17, 
    1.977246e-17, 1.994795e-17, 1.963249e-17, 1.976926e-17, 1.952144e-17, 
    1.954808e-17, 1.95964e-17, 1.970709e-17, 1.964721e-17, 1.971719e-17, 
    1.956282e-17, 1.948298e-17, 1.94622e-17, 1.942414e-17, 1.946308e-17, 
    1.945987e-17, 1.949761e-17, 1.948547e-17, 1.957619e-17, 1.952744e-17, 
    1.966598e-17, 1.971661e-17, 1.985961e-17, 1.994744e-17, 2.003673e-17, 
    2.007623e-17, 2.008825e-17, 2.009328e-17,
  8.070593e-22, 8.106384e-22, 8.099411e-22, 8.128338e-22, 8.112271e-22, 
    8.131231e-22, 8.077826e-22, 8.107822e-22, 8.088658e-22, 8.073788e-22, 
    8.184934e-22, 8.129624e-22, 8.245345e-22, 8.207946e-22, 8.302028e-22, 
    8.239539e-22, 8.314643e-22, 8.300179e-22, 8.343854e-22, 8.331175e-22, 
    8.388552e-22, 8.349792e-22, 8.418383e-22, 8.379266e-22, 8.385397e-22, 
    8.348521e-22, 8.140647e-22, 8.177802e-22, 8.138457e-22, 8.143748e-22, 
    8.141365e-22, 8.112617e-22, 8.098172e-22, 8.067833e-22, 8.07333e-22, 
    8.0956e-22, 8.146127e-22, 8.128934e-22, 8.172214e-22, 8.171234e-22, 
    8.221681e-22, 8.198667e-22, 8.28506e-22, 8.260406e-22, 8.331694e-22, 
    8.313749e-22, 8.330858e-22, 8.325664e-22, 8.330926e-22, 8.304611e-22, 
    8.315884e-22, 8.29273e-22, 8.20295e-22, 8.229227e-22, 8.152784e-22, 
    8.108564e-22, 8.079148e-22, 8.058332e-22, 8.061273e-22, 8.06689e-22, 
    8.095731e-22, 8.122852e-22, 8.143557e-22, 8.157426e-22, 8.171094e-22, 
    8.214313e-22, 8.237649e-22, 8.29007e-22, 8.280563e-22, 8.296642e-22, 
    8.311963e-22, 8.33779e-22, 8.333506e-22, 8.345145e-22, 8.296191e-22, 
    8.328556e-22, 8.275158e-22, 8.289754e-22, 8.17495e-22, 8.133564e-22, 
    8.116118e-22, 8.100756e-22, 8.063538e-22, 8.08924e-22, 8.079107e-22, 
    8.103194e-22, 8.118534e-22, 8.11094e-22, 8.157805e-22, 8.139577e-22, 
    8.239033e-22, 8.19508e-22, 8.310176e-22, 8.282511e-22, 8.316807e-22, 
    8.299292e-22, 8.329323e-22, 8.302293e-22, 8.349507e-22, 8.360059e-22, 
    8.352851e-22, 8.380507e-22, 8.300799e-22, 8.330872e-22, 8.110733e-22, 
    8.111973e-22, 8.117731e-22, 8.092435e-22, 8.090881e-22, 8.067689e-22, 
    8.088311e-22, 8.097111e-22, 8.119412e-22, 8.132641e-22, 8.145216e-22, 
    8.17289e-22, 8.205068e-22, 8.25112e-22, 8.284305e-22, 8.306587e-22, 
    8.292911e-22, 8.304986e-22, 8.291494e-22, 8.285167e-22, 8.356115e-22, 
    8.315998e-22, 8.376527e-22, 8.373131e-22, 8.34543e-22, 8.373513e-22, 
    8.11284e-22, 8.105715e-22, 8.081039e-22, 8.100347e-22, 8.065163e-22, 
    8.084867e-22, 8.096215e-22, 8.139988e-22, 8.149585e-22, 8.158531e-22, 
    8.17618e-22, 8.199836e-22, 8.2421e-22, 8.279066e-22, 8.312849e-22, 
    8.310369e-22, 8.311243e-22, 8.318812e-22, 8.300088e-22, 8.321886e-22, 
    8.325561e-22, 8.315976e-22, 8.372677e-22, 8.356269e-22, 8.373059e-22, 
    8.36237e-22, 8.108027e-22, 8.120014e-22, 8.113538e-22, 8.125725e-22, 
    8.117149e-22, 8.155349e-22, 8.166816e-22, 8.222713e-22, 8.199376e-22, 
    8.236591e-22, 8.203101e-22, 8.208967e-22, 8.237872e-22, 8.204878e-22, 
    8.277053e-22, 8.228089e-22, 8.319106e-22, 8.270166e-22, 8.32218e-22, 
    8.312703e-22, 8.328382e-22, 8.342629e-22, 8.360881e-22, 8.394644e-22, 
    8.386814e-22, 8.415057e-22, 8.137884e-22, 8.153469e-22, 8.15207e-22, 
    8.168374e-22, 8.180535e-22, 8.207937e-22, 8.252649e-22, 8.235801e-22, 
    8.266712e-22, 8.272933e-22, 8.22596e-22, 8.254813e-22, 8.163886e-22, 
    8.177912e-22, 8.16954e-22, 8.139128e-22, 8.23972e-22, 8.186864e-22, 
    8.284859e-22, 8.255939e-22, 8.340563e-22, 8.298404e-22, 8.382512e-22, 
    8.419172e-22, 8.453605e-22, 8.494063e-22, 8.161951e-22, 8.151359e-22, 
    8.170306e-22, 8.197454e-22, 8.223165e-22, 8.257707e-22, 8.26123e-22, 
    8.267717e-22, 8.284496e-22, 8.298627e-22, 8.269794e-22, 8.302169e-22, 
    8.181341e-22, 8.244334e-22, 8.147379e-22, 8.175512e-22, 8.195818e-22, 
    8.186817e-22, 8.23387e-22, 8.245072e-22, 8.290667e-22, 8.267068e-22, 
    8.410143e-22, 8.345735e-22, 8.524827e-22, 8.474646e-22, 8.147665e-22, 
    8.161903e-22, 8.213186e-22, 8.188364e-22, 8.260001e-22, 8.27777e-22, 
    8.292203e-22, 8.310712e-22, 8.312692e-22, 8.323664e-22, 8.305691e-22, 
    8.322943e-22, 8.257781e-22, 8.286871e-22, 8.207154e-22, 8.226507e-22, 
    8.21757e-22, 8.20783e-22, 8.237989e-22, 8.270255e-22, 8.270901e-22, 
    8.281266e-22, 8.31058e-22, 8.260292e-22, 8.418552e-22, 8.319784e-22, 
    8.177441e-22, 8.206227e-22, 8.2103e-22, 8.199128e-22, 8.275989e-22, 
    8.248048e-22, 8.32339e-22, 8.302992e-22, 8.336413e-22, 8.319803e-22, 
    8.317362e-22, 8.296039e-22, 8.282787e-22, 8.249337e-22, 8.22215e-22, 
    8.200743e-22, 8.205673e-22, 8.229285e-22, 8.27222e-22, 8.312891e-22, 
    8.303981e-22, 8.333871e-22, 8.254774e-22, 8.287927e-22, 8.275121e-22, 
    8.30852e-22, 8.235363e-22, 8.297776e-22, 8.219457e-22, 8.226302e-22, 
    8.247494e-22, 8.290207e-22, 8.299603e-22, 8.309721e-22, 8.303469e-22, 
    8.273303e-22, 8.268346e-22, 8.246968e-22, 8.241091e-22, 8.224808e-22, 
    8.211359e-22, 8.223658e-22, 8.236591e-22, 8.273298e-22, 8.306458e-22, 
    8.342843e-22, 8.351978e-22, 8.39584e-22, 8.360187e-22, 8.419115e-22, 
    8.369096e-22, 8.45571e-22, 8.301334e-22, 8.367539e-22, 8.248444e-22, 
    8.261129e-22, 8.284139e-22, 8.336919e-22, 8.308362e-22, 8.341896e-22, 
    8.268148e-22, 8.230124e-22, 8.220244e-22, 8.20204e-22, 8.220663e-22, 
    8.219135e-22, 8.237096e-22, 8.231321e-22, 8.274517e-22, 8.2513e-22, 
    8.317312e-22, 8.341613e-22, 8.412111e-22, 8.455475e-22, 8.499634e-22, 
    8.519182e-22, 8.525131e-22, 8.527621e-22,
  1.042633e-26, 1.047912e-26, 1.046883e-26, 1.051152e-26, 1.048781e-26, 
    1.051579e-26, 1.0437e-26, 1.048123e-26, 1.045297e-26, 1.043105e-26, 
    1.059504e-26, 1.051342e-26, 1.068305e-26, 1.062871e-26, 1.076549e-26, 
    1.067461e-26, 1.078386e-26, 1.076281e-26, 1.082654e-26, 1.080795e-26, 
    1.089248e-26, 1.08353e-26, 1.093656e-26, 1.087878e-26, 1.088783e-26, 
    1.083343e-26, 1.052971e-26, 1.058461e-26, 1.052647e-26, 1.053429e-26, 
    1.053077e-26, 1.048831e-26, 1.046699e-26, 1.042227e-26, 1.043037e-26, 
    1.04632e-26, 1.05378e-26, 1.051241e-26, 1.057637e-26, 1.057493e-26, 
    1.064868e-26, 1.061515e-26, 1.074081e-26, 1.070495e-26, 1.08087e-26, 
    1.078257e-26, 1.080748e-26, 1.079992e-26, 1.080758e-26, 1.076926e-26, 
    1.078567e-26, 1.075197e-26, 1.062141e-26, 1.065964e-26, 1.054764e-26, 
    1.048232e-26, 1.043895e-26, 1.040827e-26, 1.041261e-26, 1.042088e-26, 
    1.04634e-26, 1.050343e-26, 1.053401e-26, 1.055451e-26, 1.057472e-26, 
    1.063796e-26, 1.067187e-26, 1.074809e-26, 1.073427e-26, 1.075766e-26, 
    1.077996e-26, 1.08176e-26, 1.081134e-26, 1.082844e-26, 1.075701e-26, 
    1.080413e-26, 1.072641e-26, 1.074764e-26, 1.058039e-26, 1.051925e-26, 
    1.049347e-26, 1.047081e-26, 1.041594e-26, 1.045382e-26, 1.043888e-26, 
    1.047441e-26, 1.049705e-26, 1.048584e-26, 1.055507e-26, 1.052813e-26, 
    1.067388e-26, 1.06099e-26, 1.077736e-26, 1.07371e-26, 1.078702e-26, 
    1.076152e-26, 1.080525e-26, 1.076589e-26, 1.083488e-26, 1.085044e-26, 
    1.083981e-26, 1.088062e-26, 1.076371e-26, 1.08075e-26, 1.048554e-26, 
    1.048737e-26, 1.049587e-26, 1.045854e-26, 1.045624e-26, 1.042206e-26, 
    1.045246e-26, 1.046543e-26, 1.049835e-26, 1.051788e-26, 1.053646e-26, 
    1.057737e-26, 1.06245e-26, 1.069145e-26, 1.073971e-26, 1.077214e-26, 
    1.075223e-26, 1.076981e-26, 1.075017e-26, 1.074097e-26, 1.084462e-26, 
    1.078584e-26, 1.087475e-26, 1.086974e-26, 1.082886e-26, 1.08703e-26, 
    1.048865e-26, 1.047813e-26, 1.044173e-26, 1.047021e-26, 1.041834e-26, 
    1.044738e-26, 1.046411e-26, 1.052873e-26, 1.054292e-26, 1.055614e-26, 
    1.058224e-26, 1.061686e-26, 1.067834e-26, 1.073208e-26, 1.078126e-26, 
    1.077765e-26, 1.077892e-26, 1.078994e-26, 1.076268e-26, 1.079442e-26, 
    1.079976e-26, 1.078581e-26, 1.086906e-26, 1.084485e-26, 1.086963e-26, 
    1.085386e-26, 1.048155e-26, 1.049924e-26, 1.048968e-26, 1.050767e-26, 
    1.0495e-26, 1.055143e-26, 1.056838e-26, 1.065017e-26, 1.061618e-26, 
    1.067033e-26, 1.062163e-26, 1.063021e-26, 1.067218e-26, 1.062423e-26, 
    1.072915e-26, 1.065797e-26, 1.079037e-26, 1.071912e-26, 1.079484e-26, 
    1.078104e-26, 1.080388e-26, 1.082473e-26, 1.085166e-26, 1.090149e-26, 
    1.088993e-26, 1.093165e-26, 1.052563e-26, 1.054865e-26, 1.054659e-26, 
    1.057069e-26, 1.058864e-26, 1.06287e-26, 1.069367e-26, 1.066919e-26, 
    1.071412e-26, 1.072317e-26, 1.06549e-26, 1.069682e-26, 1.056405e-26, 
    1.058479e-26, 1.057242e-26, 1.052746e-26, 1.067488e-26, 1.059788e-26, 
    1.074051e-26, 1.069846e-26, 1.082169e-26, 1.076022e-26, 1.088358e-26, 
    1.093772e-26, 1.099017e-26, 1.105187e-26, 1.05612e-26, 1.054554e-26, 
    1.057355e-26, 1.061336e-26, 1.065084e-26, 1.070103e-26, 1.070615e-26, 
    1.071558e-26, 1.073999e-26, 1.076055e-26, 1.07186e-26, 1.076571e-26, 
    1.05898e-26, 1.068158e-26, 1.053965e-26, 1.058124e-26, 1.061098e-26, 
    1.059782e-26, 1.066639e-26, 1.068267e-26, 1.074896e-26, 1.071464e-26, 
    1.092437e-26, 1.08293e-26, 1.109886e-26, 1.102224e-26, 1.054008e-26, 
    1.056113e-26, 1.063634e-26, 1.060008e-26, 1.070436e-26, 1.07302e-26, 
    1.07512e-26, 1.077814e-26, 1.078103e-26, 1.0797e-26, 1.077083e-26, 
    1.079596e-26, 1.070113e-26, 1.074344e-26, 1.062756e-26, 1.065569e-26, 
    1.064272e-26, 1.062855e-26, 1.067237e-26, 1.071926e-26, 1.072021e-26, 
    1.073528e-26, 1.077791e-26, 1.070479e-26, 1.093678e-26, 1.079132e-26, 
    1.058411e-26, 1.062619e-26, 1.063216e-26, 1.061582e-26, 1.072761e-26, 
    1.068699e-26, 1.079661e-26, 1.07669e-26, 1.081558e-26, 1.079138e-26, 
    1.078783e-26, 1.075678e-26, 1.07375e-26, 1.068886e-26, 1.064936e-26, 
    1.061818e-26, 1.062539e-26, 1.065972e-26, 1.072212e-26, 1.078131e-26, 
    1.076834e-26, 1.081188e-26, 1.069677e-26, 1.074497e-26, 1.072634e-26, 
    1.077495e-26, 1.066855e-26, 1.075928e-26, 1.064546e-26, 1.06554e-26, 
    1.068618e-26, 1.074828e-26, 1.076197e-26, 1.07767e-26, 1.07676e-26, 
    1.07237e-26, 1.071649e-26, 1.068542e-26, 1.067688e-26, 1.065323e-26, 
    1.06337e-26, 1.065155e-26, 1.067034e-26, 1.07237e-26, 1.077195e-26, 
    1.082505e-26, 1.083852e-26, 1.090324e-26, 1.085061e-26, 1.093761e-26, 
    1.086373e-26, 1.099334e-26, 1.076447e-26, 1.086146e-26, 1.068757e-26, 
    1.0706e-26, 1.073946e-26, 1.08163e-26, 1.077472e-26, 1.082364e-26, 
    1.071621e-26, 1.066094e-26, 1.06466e-26, 1.062008e-26, 1.064721e-26, 
    1.064499e-26, 1.067108e-26, 1.066269e-26, 1.072547e-26, 1.069172e-26, 
    1.078775e-26, 1.082323e-26, 1.09273e-26, 1.099301e-26, 1.106039e-26, 
    1.109024e-26, 1.109934e-26, 1.110314e-26,
  4.215564e-32, 4.241236e-32, 4.236231e-32, 4.257018e-32, 4.24547e-32, 
    4.259101e-32, 4.22075e-32, 4.242264e-32, 4.228516e-32, 4.217859e-32, 
    4.2982e-32, 4.257945e-32, 4.341849e-32, 4.314938e-32, 4.382775e-32, 
    4.337663e-32, 4.391912e-32, 4.381449e-32, 4.413113e-32, 4.403908e-32, 
    4.445625e-32, 4.417428e-32, 4.46741e-32, 4.438868e-32, 4.443331e-32, 
    4.416504e-32, 4.265887e-32, 4.293011e-32, 4.264309e-32, 4.268117e-32, 
    4.266404e-32, 4.245715e-32, 4.235331e-32, 4.213594e-32, 4.217531e-32, 
    4.233492e-32, 4.26983e-32, 4.257455e-32, 4.288891e-32, 4.288163e-32, 
    4.324829e-32, 4.3082e-32, 4.370516e-32, 4.35272e-32, 4.404285e-32, 
    4.391275e-32, 4.403676e-32, 4.399911e-32, 4.403726e-32, 4.384656e-32, 
    4.392819e-32, 4.376062e-32, 4.311308e-32, 4.330253e-32, 4.274632e-32, 
    4.242787e-32, 4.221695e-32, 4.206793e-32, 4.208897e-32, 4.212915e-32, 
    4.233586e-32, 4.253079e-32, 4.267987e-32, 4.277986e-32, 4.288059e-32, 
    4.319512e-32, 4.336307e-32, 4.374131e-32, 4.367269e-32, 4.378885e-32, 
    4.389981e-32, 4.408704e-32, 4.405598e-32, 4.414047e-32, 4.378566e-32, 
    4.402002e-32, 4.363369e-32, 4.373911e-32, 4.290887e-32, 4.260788e-32, 
    4.248219e-32, 4.237195e-32, 4.210517e-32, 4.228929e-32, 4.221665e-32, 
    4.23895e-32, 4.249972e-32, 4.244516e-32, 4.278259e-32, 4.265118e-32, 
    4.337304e-32, 4.305589e-32, 4.388686e-32, 4.368676e-32, 4.393491e-32, 
    4.380811e-32, 4.40256e-32, 4.382982e-32, 4.417218e-32, 4.424887e-32, 
    4.419647e-32, 4.43978e-32, 4.3819e-32, 4.403683e-32, 4.244366e-32, 
    4.245256e-32, 4.249397e-32, 4.23122e-32, 4.230107e-32, 4.21349e-32, 
    4.228268e-32, 4.234578e-32, 4.250607e-32, 4.260123e-32, 4.269179e-32, 
    4.28939e-32, 4.312842e-32, 4.346016e-32, 4.369971e-32, 4.38609e-32, 
    4.376196e-32, 4.384931e-32, 4.37517e-32, 4.370598e-32, 4.422017e-32, 
    4.392899e-32, 4.43688e-32, 4.434407e-32, 4.414252e-32, 4.434686e-32, 
    4.24588e-32, 4.240762e-32, 4.223052e-32, 4.236907e-32, 4.211682e-32, 
    4.225795e-32, 4.233931e-32, 4.265406e-32, 4.272331e-32, 4.27878e-32, 
    4.291839e-32, 4.309048e-32, 4.339519e-32, 4.366182e-32, 4.390625e-32, 
    4.388829e-32, 4.389462e-32, 4.394942e-32, 4.381385e-32, 4.397171e-32, 
    4.399831e-32, 4.392888e-32, 4.434077e-32, 4.422137e-32, 4.434355e-32, 
    4.426576e-32, 4.242423e-32, 4.251037e-32, 4.246382e-32, 4.255143e-32, 
    4.248974e-32, 4.276476e-32, 4.284862e-32, 4.325561e-32, 4.308712e-32, 
    4.335551e-32, 4.311421e-32, 4.31568e-32, 4.336457e-32, 4.312714e-32, 
    4.364721e-32, 4.329423e-32, 4.395156e-32, 4.35974e-32, 4.397384e-32, 
    4.390519e-32, 4.401883e-32, 4.41222e-32, 4.425491e-32, 4.450079e-32, 
    4.444373e-32, 4.464986e-32, 4.263899e-32, 4.275125e-32, 4.274124e-32, 
    4.286034e-32, 4.295039e-32, 4.314936e-32, 4.347123e-32, 4.334991e-32, 
    4.35727e-32, 4.361758e-32, 4.327911e-32, 4.34868e-32, 4.282693e-32, 
    4.293115e-32, 4.286899e-32, 4.26479e-32, 4.337801e-32, 4.299621e-32, 
    4.37037e-32, 4.349497e-32, 4.410718e-32, 4.380158e-32, 4.441237e-32, 
    4.467976e-32, 4.494206e-32, 4.5251e-32, 4.281259e-32, 4.273611e-32, 
    4.287472e-32, 4.307309e-32, 4.325897e-32, 4.350771e-32, 4.353315e-32, 
    4.357993e-32, 4.370112e-32, 4.38033e-32, 4.359484e-32, 4.382892e-32, 
    4.295598e-32, 4.341128e-32, 4.270737e-32, 4.291328e-32, 4.306125e-32, 
    4.299596e-32, 4.333603e-32, 4.341668e-32, 4.374564e-32, 4.357528e-32, 
    4.461376e-32, 4.414465e-32, 4.549081e-32, 4.510255e-32, 4.270948e-32, 
    4.281226e-32, 4.318719e-32, 4.300719e-32, 4.352428e-32, 4.36525e-32, 
    4.375684e-32, 4.389072e-32, 4.39051e-32, 4.398457e-32, 4.385441e-32, 
    4.397938e-32, 4.350823e-32, 4.371827e-32, 4.31437e-32, 4.3283e-32, 
    4.321879e-32, 4.31486e-32, 4.336567e-32, 4.359815e-32, 4.360293e-32, 
    4.367772e-32, 4.388936e-32, 4.352639e-32, 4.467496e-32, 4.395609e-32, 
    4.292779e-32, 4.31368e-32, 4.316651e-32, 4.308538e-32, 4.363964e-32, 
    4.343809e-32, 4.398261e-32, 4.383487e-32, 4.407709e-32, 4.395661e-32, 
    4.393892e-32, 4.378457e-32, 4.368875e-32, 4.344735e-32, 4.325165e-32, 
    4.309711e-32, 4.313292e-32, 4.330297e-32, 4.361235e-32, 4.390649e-32, 
    4.384195e-32, 4.405864e-32, 4.348659e-32, 4.372584e-32, 4.363332e-32, 
    4.387487e-32, 4.334673e-32, 4.379676e-32, 4.323235e-32, 4.328157e-32, 
    4.343409e-32, 4.374225e-32, 4.381036e-32, 4.388353e-32, 4.383833e-32, 
    4.362019e-32, 4.358445e-32, 4.343033e-32, 4.338795e-32, 4.327084e-32, 
    4.317416e-32, 4.326253e-32, 4.335553e-32, 4.362021e-32, 4.385991e-32, 
    4.412373e-32, 4.419017e-32, 4.450931e-32, 4.424965e-32, 4.467905e-32, 
    4.431419e-32, 4.495774e-32, 4.382265e-32, 4.430309e-32, 4.344098e-32, 
    4.353243e-32, 4.369841e-32, 4.408059e-32, 4.387373e-32, 4.411678e-32, 
    4.358304e-32, 4.330894e-32, 4.323801e-32, 4.310651e-32, 4.324102e-32, 
    4.323004e-32, 4.335926e-32, 4.331769e-32, 4.362901e-32, 4.346156e-32, 
    4.393853e-32, 4.411475e-32, 4.462829e-32, 4.495618e-32, 4.529384e-32, 
    4.544642e-32, 4.549328e-32, 4.551289e-32,
  5.564568e-38, 5.610666e-38, 5.601667e-38, 5.639097e-38, 5.618292e-38, 
    5.642856e-38, 5.57387e-38, 5.612513e-38, 5.587805e-38, 5.568687e-38, 
    5.713715e-38, 5.640771e-38, 5.792827e-38, 5.744045e-38, 5.869254e-38, 
    5.785219e-38, 5.886477e-38, 5.86677e-38, 5.926424e-38, 5.909142e-38, 
    5.987292e-38, 5.934484e-38, 6.028307e-38, 5.974618e-38, 5.98299e-38, 
    5.932756e-38, 5.655115e-38, 5.704327e-38, 5.652263e-38, 5.65914e-38, 
    5.656048e-38, 5.618728e-38, 5.600038e-38, 5.561046e-38, 5.568099e-38, 
    5.59674e-38, 5.662235e-38, 5.639893e-38, 5.696843e-38, 5.695515e-38, 
    5.761958e-38, 5.73184e-38, 5.84621e-38, 5.81284e-38, 5.909854e-38, 
    5.885285e-38, 5.908702e-38, 5.901587e-38, 5.908794e-38, 5.872808e-38, 
    5.888197e-38, 5.856637e-38, 5.737469e-38, 5.771787e-38, 5.670923e-38, 
    5.613444e-38, 5.575563e-38, 5.548868e-38, 5.552633e-38, 5.559824e-38, 
    5.596908e-38, 5.632001e-38, 5.658913e-38, 5.676997e-38, 5.695324e-38, 
    5.752309e-38, 5.782762e-38, 5.852997e-38, 5.840116e-38, 5.86194e-38, 
    5.882847e-38, 5.918192e-38, 5.912335e-38, 5.928162e-38, 5.861348e-38, 
    5.905531e-38, 5.832799e-38, 5.852591e-38, 5.700447e-38, 5.645907e-38, 
    5.623226e-38, 5.603398e-38, 5.555532e-38, 5.588544e-38, 5.575507e-38, 
    5.606561e-38, 5.626402e-38, 5.616576e-38, 5.677492e-38, 5.653727e-38, 
    5.784574e-38, 5.727109e-38, 5.880404e-38, 5.842755e-38, 5.889466e-38, 
    5.865573e-38, 5.906587e-38, 5.86966e-38, 5.934089e-38, 5.948423e-38, 
    5.938625e-38, 5.976336e-38, 5.867623e-38, 5.908709e-38, 5.616304e-38, 
    5.617906e-38, 5.625366e-38, 5.592658e-38, 5.59066e-38, 5.560857e-38, 
    5.58736e-38, 5.598694e-38, 5.627548e-38, 5.644707e-38, 5.661065e-38, 
    5.697749e-38, 5.740243e-38, 5.800404e-38, 5.845189e-38, 5.875514e-38, 
    5.856892e-38, 5.87333e-38, 5.854961e-38, 5.84637e-38, 5.943053e-38, 
    5.888345e-38, 5.970895e-38, 5.966261e-38, 5.928544e-38, 5.966783e-38, 
    5.61903e-38, 5.60982e-38, 5.577997e-38, 5.602885e-38, 5.557621e-38, 
    5.582918e-38, 5.597525e-38, 5.654239e-38, 5.666765e-38, 5.678432e-38, 
    5.702221e-38, 5.733377e-38, 5.788601e-38, 5.83807e-38, 5.884062e-38, 
    5.880677e-38, 5.881869e-38, 5.892204e-38, 5.866653e-38, 5.896411e-38, 
    5.90143e-38, 5.888329e-38, 5.965641e-38, 5.943286e-38, 5.966163e-38, 
    5.951592e-38, 5.61281e-38, 5.628321e-38, 5.619936e-38, 5.635721e-38, 
    5.624601e-38, 5.674253e-38, 5.689481e-38, 5.763275e-38, 5.732766e-38, 
    5.781396e-38, 5.737674e-38, 5.745392e-38, 5.783024e-38, 5.74002e-38, 
    5.83532e-38, 5.770271e-38, 5.892606e-38, 5.825968e-38, 5.896814e-38, 
    5.883862e-38, 5.905314e-38, 5.924752e-38, 5.94956e-38, 5.995673e-38, 
    5.984955e-38, 6.023742e-38, 5.651525e-38, 5.671813e-38, 5.670009e-38, 
    5.691629e-38, 5.708033e-38, 5.744047e-38, 5.802422e-38, 5.780388e-38, 
    5.821363e-38, 5.829773e-38, 5.767549e-38, 5.80527e-38, 5.685535e-38, 
    5.704537e-38, 5.693204e-38, 5.653131e-38, 5.785478e-38, 5.716307e-38, 
    5.845937e-38, 5.806804e-38, 5.921948e-38, 5.864331e-38, 5.979068e-38, 
    6.029364e-38, 6.078378e-38, 6.137016e-38, 5.682924e-38, 5.669081e-38, 
    5.694255e-38, 5.730218e-38, 5.763894e-38, 5.809185e-38, 5.813953e-38, 
    5.822713e-38, 5.845457e-38, 5.864666e-38, 5.825502e-38, 5.869492e-38, 
    5.709018e-38, 5.791522e-38, 5.663879e-38, 5.701273e-38, 5.728078e-38, 
    5.716269e-38, 5.777871e-38, 5.792512e-38, 5.853814e-38, 5.821845e-38, 
    6.016918e-38, 5.928934e-38, 6.18365e-38, 6.108451e-38, 5.664264e-38, 
    5.682868e-38, 5.75089e-38, 5.718302e-38, 5.812293e-38, 5.836323e-38, 
    5.855929e-38, 5.881127e-38, 5.883844e-38, 5.898838e-38, 5.874292e-38, 
    5.897861e-38, 5.809285e-38, 5.848675e-38, 5.743022e-38, 5.76825e-38, 
    5.756622e-38, 5.743911e-38, 5.78325e-38, 5.82612e-38, 5.827028e-38, 
    5.841054e-38, 5.88083e-38, 5.812687e-38, 6.028431e-38, 5.893425e-38, 
    5.703938e-38, 5.741757e-38, 5.747154e-38, 5.732455e-38, 5.83391e-38, 
    5.796399e-38, 5.898469e-38, 5.870612e-38, 5.916329e-38, 5.893562e-38, 
    5.890222e-38, 5.861143e-38, 5.843129e-38, 5.79808e-38, 5.762568e-38, 
    5.734581e-38, 5.741069e-38, 5.771867e-38, 5.828785e-38, 5.884101e-38, 
    5.871936e-38, 5.912839e-38, 5.805238e-38, 5.850094e-38, 5.832718e-38, 
    5.878145e-38, 5.779809e-38, 5.863396e-38, 5.759078e-38, 5.767994e-38, 
    5.795673e-38, 5.853168e-38, 5.865996e-38, 5.879773e-38, 5.871262e-38, 
    5.830258e-38, 5.82356e-38, 5.794992e-38, 5.78729e-38, 5.76605e-38, 
    5.748542e-38, 5.764542e-38, 5.781403e-38, 5.830265e-38, 5.87532e-38, 
    5.925036e-38, 5.937452e-38, 5.997254e-38, 5.948555e-38, 6.0292e-38, 
    5.960609e-38, 6.081278e-38, 5.868287e-38, 5.958555e-38, 5.796927e-38, 
    5.813819e-38, 5.844935e-38, 5.916974e-38, 5.87793e-38, 5.92373e-38, 
    5.823296e-38, 5.772946e-38, 5.7601e-38, 5.736282e-38, 5.760647e-38, 
    5.758658e-38, 5.782085e-38, 5.774544e-38, 5.831917e-38, 5.800668e-38, 
    5.890145e-38, 5.923354e-38, 6.019673e-38, 6.081006e-38, 6.145331e-38, 
    6.174998e-38, 6.184138e-38, 6.187965e-38,
  2.662467e-44, 2.802597e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.662467e-44, 2.802597e-44, 2.662467e-44, 2.662467e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 
    2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.942727e-44, 2.802597e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.802597e-44, 2.802597e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.942727e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.942727e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.942727e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 3.082857e-44, 3.082857e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 3.082857e-44, 3.082857e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.802597e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 
    2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.802597e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 3.082857e-44, 2.942727e-44, 2.942727e-44, 2.802597e-44, 
    2.802597e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 2.942727e-44, 
    2.942727e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44, 2.942727e-44, 2.802597e-44, 
    2.942727e-44, 2.942727e-44, 2.942727e-44, 3.082857e-44, 3.082857e-44, 
    3.082857e-44, 3.082857e-44, 3.082857e-44,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_CH4_UNSAT =
  5.57972e-06, 5.304598e-06, 5.357845e-06, 5.137766e-06, 5.259585e-06, 
    5.115869e-06, 5.52371e-06, 5.293731e-06, 5.4403e-06, 5.554844e-06, 
    4.717595e-06, 5.128004e-06, 4.302484e-06, 4.555926e-06, 3.92762e-06, 
    4.341587e-06, 3.846678e-06, 3.939278e-06, 3.663366e-06, 3.741562e-06, 
    3.398038e-06, 3.627515e-06, 3.226016e-06, 3.452231e-06, 3.416356e-06, 
    3.635196e-06, 5.044691e-06, 4.768156e-06, 5.061202e-06, 5.021475e-06, 
    5.039296e-06, 5.257054e-06, 5.367616e-06, 5.600885e-06, 5.558384e-06, 
    5.387135e-06, 5.003639e-06, 5.133046e-06, 4.808671e-06, 4.815931e-06, 
    4.461968e-06, 4.620523e-06, 4.037266e-06, 4.199074e-06, 3.738284e-06, 
    3.852168e-06, 3.743598e-06, 3.776387e-06, 3.743172e-06, 3.910761e-06, 
    3.83859e-06, 3.987396e-06, 4.590688e-06, 4.41087e-06, 4.953641e-06, 
    5.288342e-06, 5.513574e-06, 5.674591e-06, 5.651771e-06, 5.608314e-06, 
    5.386137e-06, 5.179125e-06, 5.022709e-06, 4.918783e-06, 4.816975e-06, 
    4.512624e-06, 4.354189e-06, 4.004827e-06, 4.066543e-06, 3.96222e-06, 
    3.863576e-06, 3.700216e-06, 3.726904e-06, 3.655653e-06, 3.964973e-06, 
    3.758234e-06, 4.101852e-06, 4.006698e-06, 4.789323e-06, 5.098054e-06, 
    5.23073e-06, 5.347597e-06, 5.634236e-06, 5.435938e-06, 5.513929e-06, 
    5.328807e-06, 5.211923e-06, 5.269658e-06, 4.915949e-06, 5.052704e-06, 
    4.344858e-06, 4.645752e-06, 3.87503e-06, 4.053848e-06, 3.832648e-06, 
    3.944916e-06, 3.753352e-06, 3.925586e-06, 3.629292e-06, 3.56608e-06, 
    3.609223e-06, 3.444791e-06, 3.935222e-06, 3.743592e-06, 5.271274e-06, 
    5.261847e-06, 5.217987e-06, 5.411421e-06, 5.423311e-06, 5.602047e-06, 
    5.442954e-06, 5.375501e-06, 5.205173e-06, 5.105038e-06, 5.010317e-06, 
    4.803753e-06, 4.576054e-06, 4.263706e-06, 4.042161e-06, 3.89798e-06, 
    3.986154e-06, 3.908267e-06, 3.995372e-06, 4.036457e-06, 3.589703e-06, 
    3.837915e-06, 3.468227e-06, 3.488254e-06, 3.653963e-06, 3.485995e-06, 
    5.25523e-06, 5.30952e-06, 5.498964e-06, 5.35058e-06, 5.621585e-06, 
    5.469524e-06, 5.38249e-06, 5.049818e-06, 4.977469e-06, 4.910609e-06, 
    4.779323e-06, 4.612364e-06, 4.324089e-06, 4.076451e-06, 3.857871e-06, 
    3.873726e-06, 3.86814e-06, 3.819906e-06, 3.939819e-06, 3.800364e-06, 
    3.777152e-06, 3.837954e-06, 3.49094e-06, 3.588622e-06, 3.488681e-06, 
    3.552128e-06, 5.29186e-06, 5.200665e-06, 5.249894e-06, 5.15741e-06, 
    5.222518e-06, 4.9346e-06, 4.849132e-06, 4.455183e-06, 4.615629e-06, 
    4.361188e-06, 4.589575e-06, 4.548821e-06, 4.352937e-06, 4.57714e-06, 
    4.089787e-06, 4.418833e-06, 3.818036e-06, 4.135183e-06, 3.798496e-06, 
    3.858805e-06, 3.759171e-06, 3.670854e-06, 3.561047e-06, 3.362361e-06, 
    3.407903e-06, 3.244832e-06, 5.065449e-06, 4.948547e-06, 4.958825e-06, 
    4.837228e-06, 4.74785e-06, 4.555872e-06, 4.253386e-06, 4.366312e-06, 
    4.15741e-06, 4.11654e-06, 4.432807e-06, 4.239027e-06, 4.870737e-06, 
    4.766819e-06, 4.828625e-06, 5.056192e-06, 4.340179e-06, 4.703499e-06, 
    4.038579e-06, 4.231405e-06, 3.68339e-06, 3.95089e-06, 3.433093e-06, 
    3.221739e-06, 3.028965e-06, 2.811587e-06, 4.885075e-06, 4.964151e-06, 
    4.822828e-06, 4.629233e-06, 4.451867e-06, 4.219668e-06, 4.193619e-06, 
    4.150852e-06, 4.040845e-06, 3.949218e-06, 4.137348e-06, 3.926379e-06, 
    4.742781e-06, 4.30911e-06, 4.994123e-06, 4.784621e-06, 4.640585e-06, 
    4.703622e-06, 4.379287e-06, 4.303965e-06, 4.000906e-06, 4.155056e-06, 
    3.273289e-06, 3.652295e-06, 2.652207e-06, 2.914831e-06, 4.991857e-06, 
    4.885354e-06, 4.519918e-06, 4.692728e-06, 4.201753e-06, 4.08485e-06, 
    3.990741e-06, 3.871662e-06, 3.858902e-06, 3.789127e-06, 3.903734e-06, 
    3.793633e-06, 4.219178e-06, 4.025433e-06, 4.561264e-06, 4.429198e-06, 
    4.489798e-06, 4.556573e-06, 4.351542e-06, 4.134357e-06, 4.12985e-06, 
    4.062073e-06, 3.873361e-06, 4.19982e-06, 3.225761e-06, 3.814517e-06, 
    4.769954e-06, 4.568091e-06, 4.539509e-06, 4.617231e-06, 4.096515e-06, 
    4.284103e-06, 3.790825e-06, 3.921088e-06, 3.708608e-06, 3.813584e-06, 
    3.82913e-06, 3.965935e-06, 4.052051e-06, 4.275533e-06, 4.458791e-06, 
    4.605936e-06, 4.571585e-06, 4.410437e-06, 4.121397e-06, 3.857737e-06, 
    3.914907e-06, 3.724584e-06, 4.239124e-06, 4.018679e-06, 4.102322e-06, 
    3.885629e-06, 4.369322e-06, 3.955543e-06, 4.476952e-06, 4.430492e-06, 
    4.287814e-06, 4.004052e-06, 3.942919e-06, 3.878013e-06, 3.918018e-06, 
    4.114238e-06, 4.146741e-06, 4.291268e-06, 4.330805e-06, 4.440596e-06, 
    4.532172e-06, 4.448472e-06, 4.361127e-06, 4.114165e-06, 3.898942e-06, 
    3.6696e-06, 3.614379e-06, 3.355818e-06, 3.565611e-06, 3.222606e-06, 
    3.513153e-06, 3.018039e-06, 3.932254e-06, 3.52192e-06, 4.281368e-06, 
    4.194271e-06, 4.043459e-06, 3.705782e-06, 3.886638e-06, 3.675496e-06, 
    4.148018e-06, 4.404899e-06, 4.471621e-06, 4.596942e-06, 4.468769e-06, 
    4.47915e-06, 4.357539e-06, 4.396498e-06, 4.106158e-06, 4.262282e-06, 
    3.829515e-06, 3.67715e-06, 3.261733e-06, 3.01895e-06, 2.782044e-06, 
    2.680908e-06, 2.650563e-06, 2.637937e-06,
  8.252538e-06, 8.083487e-06, 8.116155e-06, 7.981281e-06, 8.055884e-06, 
    7.967883e-06, 8.21807e-06, 8.076826e-06, 8.166791e-06, 8.237223e-06, 
    7.724962e-06, 7.975306e-06, 7.473346e-06, 7.626751e-06, 6.964633e-06, 
    7.496975e-06, 6.92643e-06, 6.970137e-06, 6.840277e-06, 6.876962e-06, 
    6.716518e-06, 6.823489e-06, 6.636868e-06, 6.741703e-06, 6.725024e-06, 
    6.827085e-06, 7.924356e-06, 7.755722e-06, 7.934449e-06, 7.910175e-06, 
    7.92106e-06, 8.054335e-06, 8.122161e-06, 8.265562e-06, 8.239402e-06, 
    8.13414e-06, 7.899281e-06, 7.978387e-06, 7.780362e-06, 7.784784e-06, 
    7.569799e-06, 7.665951e-06, 7.016533e-06, 7.093465e-06, 6.875423e-06, 
    6.929013e-06, 6.87792e-06, 6.89333e-06, 6.877719e-06, 6.956662e-06, 
    6.922614e-06, 6.992901e-06, 7.647842e-06, 7.538866e-06, 7.868752e-06, 
    8.07353e-06, 8.211837e-06, 8.310967e-06, 8.296905e-06, 8.270141e-06, 
    8.133527e-06, 8.006591e-06, 7.910923e-06, 7.847479e-06, 7.785421e-06, 
    7.600509e-06, 7.504588e-06, 7.001161e-06, 7.030423e-06, 6.980989e-06, 
    6.934391e-06, 6.857555e-06, 6.870079e-06, 6.836666e-06, 6.982288e-06, 
    6.884799e-06, 7.047191e-06, 7.002043e-06, 7.768609e-06, 7.956981e-06, 
    8.038213e-06, 8.109868e-06, 8.286104e-06, 8.164115e-06, 8.212057e-06, 
    8.098333e-06, 8.026678e-06, 8.062057e-06, 7.84575e-06, 7.929253e-06, 
    7.498947e-06, 7.681278e-06, 6.939794e-06, 7.024398e-06, 6.919813e-06, 
    6.9728e-06, 6.882504e-06, 6.963664e-06, 6.824323e-06, 6.794772e-06, 
    6.814934e-06, 6.738238e-06, 6.968218e-06, 6.877919e-06, 8.063049e-06, 
    8.05727e-06, 8.030392e-06, 8.149053e-06, 8.156356e-06, 8.26628e-06, 
    8.168421e-06, 8.126995e-06, 8.022541e-06, 7.961252e-06, 7.903354e-06, 
    7.77737e-06, 7.638965e-06, 7.449931e-06, 7.018854e-06, 6.950624e-06, 
    6.992311e-06, 6.955482e-06, 6.996677e-06, 7.016147e-06, 6.80581e-06, 
    6.922297e-06, 6.749143e-06, 6.758469e-06, 6.835876e-06, 6.757416e-06, 
    8.053215e-06, 8.0865e-06, 8.202851e-06, 8.111693e-06, 8.278311e-06, 
    8.184753e-06, 8.131289e-06, 7.927495e-06, 7.883293e-06, 7.842495e-06, 
    7.762495e-06, 7.660998e-06, 7.486392e-06, 7.035129e-06, 6.9317e-06, 
    6.939177e-06, 6.936543e-06, 6.913811e-06, 6.970391e-06, 6.904611e-06, 
    6.893693e-06, 6.922313e-06, 6.75972e-06, 6.8053e-06, 6.758667e-06, 
    6.788254e-06, 8.075669e-06, 8.019781e-06, 8.049943e-06, 7.993299e-06, 
    8.03317e-06, 7.857137e-06, 7.805023e-06, 7.565697e-06, 7.662981e-06, 
    7.508816e-06, 7.647164e-06, 7.622442e-06, 7.503839e-06, 7.639617e-06, 
    7.041467e-06, 7.543693e-06, 6.912931e-06, 7.063053e-06, 6.903732e-06, 
    6.93214e-06, 6.885236e-06, 6.843788e-06, 6.792419e-06, 6.699955e-06, 
    6.721093e-06, 6.645553e-06, 7.937043e-06, 7.865644e-06, 7.871911e-06, 
    7.797759e-06, 7.743343e-06, 7.626715e-06, 7.443699e-06, 7.511908e-06, 
    7.073617e-06, 7.054175e-06, 7.552138e-06, 7.435039e-06, 7.818184e-06, 
    7.754894e-06, 7.79252e-06, 7.931389e-06, 7.496117e-06, 7.716375e-06, 
    7.017156e-06, 7.430438e-06, 6.849665e-06, 6.975632e-06, 6.7328e-06, 
    6.634899e-06, 6.546237e-06, 6.447074e-06, 7.826923e-06, 7.875162e-06, 
    7.788985e-06, 7.671247e-06, 7.563681e-06, 7.423361e-06, 7.090865e-06, 
    7.070497e-06, 7.018228e-06, 6.974835e-06, 7.064076e-06, 6.964038e-06, 
    7.740278e-06, 7.477343e-06, 7.893465e-06, 7.765731e-06, 7.678139e-06, 
    7.716443e-06, 7.519753e-06, 7.47423e-06, 6.999303e-06, 7.072496e-06, 
    6.658714e-06, 6.835099e-06, 6.374947e-06, 6.494063e-06, 7.892078e-06, 
    7.82709e-06, 7.604919e-06, 7.709819e-06, 7.094742e-06, 7.039117e-06, 
    6.994484e-06, 6.938207e-06, 6.932187e-06, 6.899324e-06, 6.953341e-06, 
    6.901443e-06, 7.423066e-06, 7.010921e-06, 7.629984e-06, 7.549956e-06, 
    7.586656e-06, 7.627139e-06, 7.502977e-06, 7.062654e-06, 7.060503e-06, 
    7.028304e-06, 6.939031e-06, 7.09382e-06, 6.636768e-06, 6.911294e-06, 
    7.756791e-06, 7.634137e-06, 7.616793e-06, 7.66395e-06, 7.044658e-06, 
    7.462239e-06, 6.900123e-06, 6.961538e-06, 6.861491e-06, 6.910834e-06, 
    6.918156e-06, 6.982742e-06, 7.023546e-06, 7.457067e-06, 7.567875e-06, 
    7.657092e-06, 7.636246e-06, 7.538602e-06, 7.056488e-06, 6.93164e-06, 
    6.958623e-06, 6.868989e-06, 7.435093e-06, 7.007723e-06, 7.04742e-06, 
    6.944796e-06, 7.51373e-06, 6.977848e-06, 7.578873e-06, 7.550737e-06, 
    7.464479e-06, 7.000797e-06, 6.971857e-06, 6.941204e-06, 6.960087e-06, 
    7.053084e-06, 7.068541e-06, 7.466563e-06, 7.490448e-06, 7.556853e-06, 
    7.612341e-06, 7.561624e-06, 7.508777e-06, 7.053046e-06, 6.951082e-06, 
    6.843201e-06, 6.817344e-06, 6.696931e-06, 6.794561e-06, 6.635314e-06, 
    6.770098e-06, 6.541247e-06, 6.966828e-06, 6.774173e-06, 7.460585e-06, 
    7.091175e-06, 7.019476e-06, 6.860173e-06, 6.945271e-06, 6.845969e-06, 
    7.069149e-06, 7.535256e-06, 7.575643e-06, 7.651634e-06, 7.573916e-06, 
    7.580205e-06, 7.506602e-06, 7.530163e-06, 7.04924e-06, 7.449064e-06, 
    6.918339e-06, 6.846743e-06, 6.653364e-06, 6.541655e-06, 6.433658e-06, 
    6.387893e-06, 6.374203e-06, 6.368513e-06,
  9.62226e-06, 9.637781e-06, 9.634949e-06, 9.646082e-06, 9.640107e-06, 
    9.647105e-06, 9.625596e-06, 9.638346e-06, 9.630399e-06, 9.623754e-06, 
    9.662808e-06, 9.64654e-06, 9.672562e-06, 9.667482e-06, 1.000894e-05, 
    9.671965e-06, 9.994018e-06, 1.001107e-05, 9.959294e-06, 9.974269e-06, 
    9.906511e-06, 9.952344e-06, 9.870474e-06, 9.917555e-06, 9.91026e-06, 
    9.953837e-06, 9.650324e-06, 9.661136e-06, 9.649592e-06, 9.651335e-06, 
    9.65056e-06, 9.640235e-06, 9.634418e-06, 9.620979e-06, 9.623543e-06, 
    9.633355e-06, 9.6521e-06, 9.646305e-06, 9.659732e-06, 9.659473e-06, 
    9.669697e-06, 9.665744e-06, 1.002879e-05, 1.005736e-05, 9.973646e-06, 
    9.995038e-06, 9.974656e-06, 9.980859e-06, 9.974575e-06, 1.000586e-05, 
    9.992514e-06, 1.001982e-05, 9.666568e-06, 9.67074e-06, 9.654187e-06, 
    9.638625e-06, 9.62619e-06, 9.616418e-06, 9.617846e-06, 9.620525e-06, 
    9.63341e-06, 9.644108e-06, 9.651283e-06, 9.65559e-06, 9.659436e-06, 
    9.668545e-06, 9.671759e-06, 1.002296e-05, 1.003402e-05, 1.001525e-05, 
    9.997154e-06, 9.966382e-06, 9.971481e-06, 9.957804e-06, 1.001575e-05, 
    9.97743e-06, 1.004029e-05, 1.00233e-05, 9.660405e-06, 9.647928e-06, 
    9.641562e-06, 9.635501e-06, 9.618932e-06, 9.630644e-06, 9.626168e-06, 
    9.636506e-06, 9.642502e-06, 9.639593e-06, 9.655702e-06, 9.649971e-06, 
    9.671913e-06, 9.665018e-06, 9.999274e-06, 1.003176e-05, 9.991407e-06, 
    1.00121e-05, 9.976506e-06, 1.000857e-05, 9.95269e-06, 9.940307e-06, 
    9.948777e-06, 9.916047e-06, 1.001033e-05, 9.974654e-06, 9.63951e-06, 
    9.639993e-06, 9.642202e-06, 9.632015e-06, 9.631352e-06, 9.620908e-06, 
    9.63025e-06, 9.633992e-06, 9.642836e-06, 9.647607e-06, 9.651816e-06, 
    9.659906e-06, 9.666957e-06, 9.673082e-06, 1.002967e-05, 1.000351e-05, 
    1.001959e-05, 1.00054e-05, 1.002126e-05, 1.002865e-05, 9.944954e-06, 
    9.992388e-06, 9.920788e-06, 9.924818e-06, 9.957476e-06, 9.924365e-06, 
    9.640329e-06, 9.637524e-06, 9.627041e-06, 9.635342e-06, 9.619713e-06, 
    9.628739e-06, 9.633609e-06, 9.650096e-06, 9.653205e-06, 9.655912e-06, 
    9.66076e-06, 9.665973e-06, 9.672242e-06, 1.003579e-05, 9.996097e-06, 
    9.999033e-06, 9.998e-06, 9.989029e-06, 1.001117e-05, 9.98537e-06, 
    9.981003e-06, 9.992395e-06, 9.925358e-06, 9.944742e-06, 9.924905e-06, 
    9.937551e-06, 9.638446e-06, 9.643057e-06, 9.6406e-06, 9.645151e-06, 
    9.641975e-06, 9.654957e-06, 9.658259e-06, 9.66984e-06, 9.665881e-06, 
    9.671642e-06, 9.666599e-06, 9.667662e-06, 9.671778e-06, 9.666931e-06, 
    1.003816e-05, 9.670583e-06, 9.988679e-06, 1.004618e-05, 9.985019e-06, 
    9.99627e-06, 9.977607e-06, 9.960739e-06, 9.939314e-06, 9.899162e-06, 
    9.908533e-06, 9.874492e-06, 9.649403e-06, 9.654394e-06, 9.653976e-06, 
    9.658701e-06, 9.661826e-06, 9.667484e-06, 9.673209e-06, 9.671556e-06, 
    1.005008e-05, 1.004289e-05, 9.670308e-06, 9.673376e-06, 9.657451e-06, 
    9.661186e-06, 9.659014e-06, 9.649815e-06, 9.67199e-06, 9.663261e-06, 
    1.002903e-05, 9.673461e-06, 9.963152e-06, 1.001319e-05, 9.913671e-06, 
    9.869557e-06, 9.827168e-06, 9.776493e-06, 9.656905e-06, 9.653757e-06, 
    9.659225e-06, 9.665495e-06, 9.669912e-06, 9.673586e-06, 1.005641e-05, 
    1.004893e-05, 1.002943e-05, 1.001289e-05, 1.004656e-05, 1.000872e-05, 
    9.661988e-06, 9.672467e-06, 9.652505e-06, 9.660574e-06, 9.665168e-06, 
    9.663259e-06, 9.671328e-06, 9.672543e-06, 1.002226e-05, 1.004967e-05, 
    9.880531e-06, 9.957153e-06, 9.737092e-06, 9.800971e-06, 9.652601e-06, 
    9.656895e-06, 9.668374e-06, 9.6636e-06, 1.005782e-05, 1.003728e-05, 
    1.002042e-05, 9.998651e-06, 9.996288e-06, 9.983259e-06, 1.000456e-05, 
    9.984105e-06, 9.67359e-06, 1.002667e-05, 9.667346e-06, 9.67038e-06, 
    9.669081e-06, 9.667467e-06, 9.671806e-06, 1.004603e-05, 1.004524e-05, 
    1.003323e-05, 9.998964e-06, 1.005749e-05, 9.870418e-06, 9.98802e-06, 
    9.661082e-06, 9.667166e-06, 9.667897e-06, 9.665838e-06, 1.003935e-05, 
    9.672819e-06, 9.983578e-06, 1.000775e-05, 9.967988e-06, 9.987846e-06, 
    9.990751e-06, 1.001593e-05, 1.003144e-05, 9.672932e-06, 9.669765e-06, 
    9.666152e-06, 9.667077e-06, 9.670748e-06, 1.004375e-05, 9.996072e-06, 
    1.000662e-05, 9.971039e-06, 9.673376e-06, 1.002546e-05, 1.004038e-05, 
    1.000123e-05, 9.671503e-06, 1.001404e-05, 9.66937e-06, 9.670354e-06, 
    9.672769e-06, 1.002282e-05, 1.001174e-05, 9.999825e-06, 1.000719e-05, 
    1.004248e-05, 1.004821e-05, 9.672722e-06, 9.67214e-06, 9.670149e-06, 
    9.668079e-06, 9.669984e-06, 9.671644e-06, 1.004247e-05, 1.000368e-05, 
    9.960497e-06, 9.949785e-06, 9.897807e-06, 9.940214e-06, 9.869742e-06, 
    9.929802e-06, 9.824696e-06, 1.000979e-05, 9.931551e-06, 9.672856e-06, 
    1.005652e-05, 1.00299e-05, 9.967447e-06, 1.000142e-05, 9.961633e-06, 
    1.004843e-05, 9.670854e-06, 9.669488e-06, 9.666399e-06, 9.66955e-06, 
    9.669321e-06, 9.671706e-06, 9.671015e-06, 1.004106e-05, 9.673102e-06, 
    9.990823e-06, 9.961952e-06, 9.878085e-06, 9.824903e-06, 9.769344e-06, 
    9.744343e-06, 9.736675e-06, 9.733461e-06,
  4.406788e-06, 4.320465e-06, 4.337236e-06, 4.267702e-06, 4.306263e-06, 
    4.26075e-06, 4.389278e-06, 4.317038e-06, 4.363143e-06, 4.399015e-06, 
    4.13311e-06, 4.264604e-06, 3.997116e-06, 4.080557e-06, 3.871733e-06, 
    4.01008e-06, 3.843867e-06, 3.875731e-06, 3.779983e-06, 3.807372e-06, 
    3.685351e-06, 3.767354e-06, 3.622408e-06, 3.704909e-06, 3.691976e-06, 
    3.770064e-06, 4.238111e-06, 4.149451e-06, 4.243369e-06, 4.230712e-06, 
    4.236393e-06, 4.305463e-06, 4.340308e-06, 4.413398e-06, 4.400122e-06, 
    4.346447e-06, 4.225022e-06, 4.266205e-06, 4.162518e-06, 4.164856e-06, 
    4.049781e-06, 4.101614e-06, 3.909176e-06, 3.963835e-06, 3.806228e-06, 
    3.845764e-06, 3.808082e-06, 3.819503e-06, 3.807934e-06, 3.865946e-06, 
    3.841072e-06, 3.892188e-06, 4.091898e-06, 4.032967e-06, 4.209047e-06, 
    4.315337e-06, 4.386106e-06, 4.436381e-06, 4.42927e-06, 4.415716e-06, 
    4.346133e-06, 4.280815e-06, 4.231106e-06, 4.19789e-06, 4.165192e-06, 
    4.066394e-06, 4.014251e-06, 3.898133e-06, 3.919116e-06, 3.883586e-06, 
    3.849702e-06, 3.792916e-06, 3.802254e-06, 3.77727e-06, 3.884528e-06, 
    3.813184e-06, 3.931075e-06, 3.898772e-06, 4.156279e-06, 4.255091e-06, 
    4.297144e-06, 4.33401e-06, 4.423803e-06, 4.361774e-06, 4.386216e-06, 
    4.328094e-06, 4.291198e-06, 4.309444e-06, 4.196982e-06, 4.240664e-06, 
    4.011163e-06, 4.109816e-06, 3.853651e-06, 3.914809e-06, 3.839017e-06, 
    3.877663e-06, 3.811483e-06, 3.871036e-06, 3.767981e-06, 3.745602e-06, 
    3.760892e-06, 3.702232e-06, 3.874341e-06, 3.80808e-06, 4.309954e-06, 
    4.306977e-06, 4.293116e-06, 4.354077e-06, 4.357811e-06, 4.413761e-06, 
    4.363976e-06, 4.342789e-06, 4.289062e-06, 4.257311e-06, 4.227153e-06, 
    4.160933e-06, 4.087126e-06, 3.984227e-06, 3.910839e-06, 3.861553e-06, 
    3.891765e-06, 3.86509e-06, 3.89491e-06, 3.908901e-06, 3.753983e-06, 
    3.840838e-06, 3.710658e-06, 3.717842e-06, 3.776675e-06, 3.717032e-06, 
    4.304888e-06, 4.322017e-06, 4.381531e-06, 4.33495e-06, 4.419857e-06, 
    4.372308e-06, 4.344986e-06, 4.239744e-06, 4.216666e-06, 4.19527e-06, 
    4.153057e-06, 4.098958e-06, 4.004285e-06, 3.922475e-06, 3.847733e-06, 
    3.853202e-06, 3.851276e-06, 3.834606e-06, 3.875917e-06, 3.827832e-06, 
    3.819769e-06, 3.840853e-06, 3.718804e-06, 3.7536e-06, 3.717994e-06, 
    3.740644e-06, 4.316449e-06, 4.287635e-06, 4.303202e-06, 4.273933e-06, 
    4.294549e-06, 4.202954e-06, 4.175536e-06, 4.047551e-06, 4.100021e-06, 
    4.016566e-06, 4.091535e-06, 4.078236e-06, 4.013836e-06, 4.087481e-06, 
    3.926991e-06, 4.03559e-06, 3.833959e-06, 3.942331e-06, 3.827183e-06, 
    3.848056e-06, 3.813511e-06, 3.782615e-06, 3.743815e-06, 3.672408e-06, 
    3.688922e-06, 3.629361e-06, 4.244721e-06, 4.207418e-06, 4.210706e-06, 
    4.17171e-06, 4.142896e-06, 4.080539e-06, 3.980791e-06, 4.018261e-06, 
    3.949825e-06, 3.936039e-06, 4.040193e-06, 3.976005e-06, 4.182478e-06, 
    4.149021e-06, 4.168941e-06, 4.241774e-06, 4.009614e-06, 4.128548e-06, 
    3.909622e-06, 3.973464e-06, 3.787017e-06, 3.879708e-06, 3.698017e-06, 
    3.620824e-06, 3.5485e-06, 3.464341e-06, 4.187081e-06, 4.212409e-06, 
    4.167076e-06, 4.104446e-06, 4.046462e-06, 3.969546e-06, 3.962003e-06, 
    3.947615e-06, 3.910393e-06, 3.879137e-06, 3.943062e-06, 3.871308e-06, 
    4.141255e-06, 3.999317e-06, 4.221984e-06, 4.154765e-06, 4.108137e-06, 
    4.128589e-06, 4.022549e-06, 3.99761e-06, 3.896797e-06, 3.949032e-06, 
    3.639841e-06, 3.776087e-06, 3.400583e-06, 3.504686e-06, 4.221261e-06, 
    4.187171e-06, 4.068784e-06, 4.12506e-06, 3.964734e-06, 3.925321e-06, 
    3.893331e-06, 3.85249e-06, 3.848089e-06, 3.82393e-06, 3.863531e-06, 
    3.825496e-06, 3.969382e-06, 3.905152e-06, 4.082301e-06, 4.039005e-06, 
    4.058917e-06, 4.080769e-06, 4.013377e-06, 3.942053e-06, 3.940534e-06, 
    3.9176e-06, 3.853072e-06, 3.964085e-06, 3.62231e-06, 3.832736e-06, 
    4.150035e-06, 4.084527e-06, 4.075193e-06, 4.100543e-06, 3.929269e-06, 
    3.991012e-06, 3.82452e-06, 3.869493e-06, 3.795855e-06, 3.832416e-06, 
    3.8378e-06, 3.884857e-06, 3.914199e-06, 3.988162e-06, 4.048738e-06, 
    4.096866e-06, 4.085669e-06, 4.032825e-06, 3.937679e-06, 3.847686e-06, 
    3.867369e-06, 3.801443e-06, 3.976038e-06, 3.902852e-06, 3.931233e-06, 
    3.857303e-06, 4.019256e-06, 3.881298e-06, 4.054702e-06, 4.039431e-06, 
    3.992246e-06, 3.897868e-06, 3.876979e-06, 3.854679e-06, 3.868439e-06, 
    3.935261e-06, 3.94623e-06, 3.993393e-06, 4.00651e-06, 4.042756e-06, 
    4.072794e-06, 4.045346e-06, 4.016546e-06, 3.935237e-06, 3.861883e-06, 
    3.782174e-06, 3.762715e-06, 3.670026e-06, 3.745434e-06, 3.621142e-06, 
    3.726744e-06, 3.544335e-06, 3.873321e-06, 3.729877e-06, 3.990103e-06, 
    3.962222e-06, 3.91128e-06, 3.794864e-06, 3.85765e-06, 3.784245e-06, 
    3.946661e-06, 4.030999e-06, 4.052952e-06, 4.093936e-06, 4.052016e-06, 
    4.055423e-06, 4.01536e-06, 4.028229e-06, 3.932531e-06, 3.983754e-06, 
    3.837933e-06, 3.784826e-06, 3.635591e-06, 3.544685e-06, 3.452666e-06, 
    3.412207e-06, 3.399916e-06, 3.39478e-06,
  4.550293e-07, 4.380055e-07, 4.412853e-07, 4.277731e-07, 4.352384e-07, 
    4.264347e-07, 4.515476e-07, 4.373369e-07, 4.463781e-07, 4.53482e-07, 
    4.022619e-07, 4.271763e-07, 3.773407e-07, 3.9253e-07, 3.550694e-07, 
    3.796794e-07, 3.502304e-07, 3.557668e-07, 3.392699e-07, 3.439463e-07, 
    3.233738e-07, 3.371252e-07, 3.130245e-07, 3.26626e-07, 3.244735e-07, 
    3.375847e-07, 4.220918e-07, 4.053142e-07, 4.230982e-07, 4.206774e-07, 
    4.21763e-07, 4.350828e-07, 4.418876e-07, 4.563474e-07, 4.537021e-07, 
    4.430923e-07, 4.195916e-07, 4.274847e-07, 4.07764e-07, 4.082032e-07, 
    3.868902e-07, 3.964141e-07, 3.616275e-07, 3.713161e-07, 3.437503e-07, 
    3.505588e-07, 3.44068e-07, 3.460284e-07, 3.440425e-07, 3.540617e-07, 
    3.49747e-07, 3.586443e-07, 3.946194e-07, 3.838275e-07, 4.165515e-07, 
    4.370052e-07, 4.509184e-07, 4.609465e-07, 4.595209e-07, 4.568101e-07, 
    4.430307e-07, 4.303039e-07, 4.207527e-07, 4.14435e-07, 4.082664e-07, 
    3.899292e-07, 3.804336e-07, 3.596867e-07, 3.633793e-07, 3.571385e-07, 
    3.512407e-07, 3.414739e-07, 3.430698e-07, 3.388085e-07, 3.573033e-07, 
    3.44943e-07, 3.654928e-07, 3.597988e-07, 4.065933e-07, 4.253469e-07, 
    4.334666e-07, 4.406535e-07, 4.584265e-07, 4.461081e-07, 4.509404e-07, 
    4.394959e-07, 4.323136e-07, 4.358573e-07, 4.142631e-07, 4.225802e-07, 
    3.798752e-07, 3.979326e-07, 3.519255e-07, 3.626197e-07, 3.493918e-07, 
    3.561039e-07, 3.446511e-07, 3.549481e-07, 3.372314e-07, 3.334479e-07, 
    3.360304e-07, 3.261798e-07, 3.555243e-07, 3.440676e-07, 4.359566e-07, 
    4.353773e-07, 4.326854e-07, 4.445923e-07, 4.453272e-07, 4.564197e-07, 
    4.465423e-07, 4.423743e-07, 4.318998e-07, 4.257733e-07, 4.199982e-07, 
    4.074665e-07, 3.937395e-07, 3.750229e-07, 3.619204e-07, 3.532976e-07, 
    3.5857e-07, 3.539126e-07, 3.591214e-07, 3.615791e-07, 3.348621e-07, 
    3.497066e-07, 3.275853e-07, 3.287859e-07, 3.387073e-07, 3.286505e-07, 
    4.34971e-07, 4.383085e-07, 4.50012e-07, 4.408375e-07, 4.576375e-07, 
    4.481872e-07, 4.428055e-07, 4.224041e-07, 4.179999e-07, 4.139389e-07, 
    4.059897e-07, 3.959232e-07, 3.786329e-07, 3.639722e-07, 3.508997e-07, 
    3.518476e-07, 3.515136e-07, 3.486301e-07, 3.557991e-07, 3.474618e-07, 
    3.460741e-07, 3.49709e-07, 3.289469e-07, 3.347975e-07, 3.288115e-07, 
    3.326126e-07, 4.372221e-07, 4.316235e-07, 4.346433e-07, 4.289747e-07, 
    4.329632e-07, 4.153949e-07, 4.102124e-07, 3.864832e-07, 3.961195e-07, 
    3.808526e-07, 3.945525e-07, 3.921031e-07, 3.803584e-07, 3.93805e-07, 
    3.647702e-07, 3.843043e-07, 3.485183e-07, 3.67488e-07, 3.473501e-07, 
    3.509556e-07, 3.449992e-07, 3.397178e-07, 3.331467e-07, 3.212311e-07, 
    3.239663e-07, 3.14159e-07, 4.233573e-07, 4.16242e-07, 4.168666e-07, 
    4.094919e-07, 4.040885e-07, 3.925268e-07, 3.744064e-07, 3.811595e-07, 
    3.688197e-07, 3.663721e-07, 3.851421e-07, 3.735485e-07, 4.115213e-07, 
    4.052339e-07, 4.089711e-07, 4.227928e-07, 3.795953e-07, 4.014121e-07, 
    3.61706e-07, 3.730933e-07, 3.404676e-07, 3.56461e-07, 3.254779e-07, 
    3.127663e-07, 3.01099e-07, 2.878165e-07, 4.123904e-07, 4.171903e-07, 
    4.086205e-07, 3.96938e-07, 3.862846e-07, 3.723923e-07, 3.709891e-07, 
    3.684268e-07, 3.618417e-07, 3.563611e-07, 3.676179e-07, 3.549955e-07, 
    4.037819e-07, 3.777371e-07, 4.190127e-07, 4.063095e-07, 3.976214e-07, 
    4.014198e-07, 3.819362e-07, 3.774296e-07, 3.594523e-07, 3.686787e-07, 
    3.158731e-07, 3.386074e-07, 2.779633e-07, 2.941445e-07, 4.18875e-07, 
    4.124074e-07, 3.903674e-07, 4.007629e-07, 3.714766e-07, 3.64475e-07, 
    3.588445e-07, 3.517241e-07, 3.509613e-07, 3.4679e-07, 3.536416e-07, 
    3.470594e-07, 3.723631e-07, 3.609196e-07, 3.928509e-07, 3.849257e-07, 
    3.885598e-07, 3.92569e-07, 3.802755e-07, 3.674388e-07, 3.671691e-07, 
    3.631117e-07, 3.518249e-07, 3.713608e-07, 3.130084e-07, 3.483072e-07, 
    4.054236e-07, 3.932608e-07, 3.915439e-07, 3.962161e-07, 3.651732e-07, 
    3.762421e-07, 3.468915e-07, 3.546792e-07, 3.419758e-07, 3.482522e-07, 
    3.491815e-07, 3.573609e-07, 3.625121e-07, 3.757298e-07, 3.866997e-07, 
    3.955365e-07, 3.934711e-07, 3.838016e-07, 3.666627e-07, 3.508916e-07, 
    3.543094e-07, 3.429311e-07, 3.735545e-07, 3.605154e-07, 3.655207e-07, 
    3.525591e-07, 3.813396e-07, 3.567386e-07, 3.877891e-07, 3.850034e-07, 
    3.764639e-07, 3.596403e-07, 3.559845e-07, 3.521037e-07, 3.544956e-07, 
    3.662342e-07, 3.681806e-07, 3.766705e-07, 3.790346e-07, 3.85609e-07, 
    3.911034e-07, 3.860811e-07, 3.808489e-07, 3.662298e-07, 3.53355e-07, 
    3.396428e-07, 3.363391e-07, 3.208376e-07, 3.334195e-07, 3.128181e-07, 
    3.302771e-07, 3.004342e-07, 3.553464e-07, 3.308028e-07, 3.760787e-07, 
    3.710282e-07, 3.619978e-07, 3.418065e-07, 3.526195e-07, 3.399953e-07, 
    3.682571e-07, 3.834697e-07, 3.874693e-07, 3.949955e-07, 3.872983e-07, 
    3.879209e-07, 3.806344e-07, 3.829668e-07, 3.657505e-07, 3.749381e-07, 
    3.492045e-07, 3.400942e-07, 3.151773e-07, 3.0049e-07, 2.859987e-07, 
    2.797463e-07, 2.778611e-07, 2.770754e-07,
  1.281292e-08, 1.207717e-08, 1.221774e-08, 1.164227e-08, 1.195902e-08, 
    1.15858e-08, 1.266122e-08, 1.204859e-08, 1.243714e-08, 1.274542e-08, 
    1.058242e-08, 1.161708e-08, 9.581544e-09, 1.018746e-08, 8.71681e-09, 
    9.673993e-09, 8.532718e-09, 8.743451e-09, 8.120851e-09, 8.295707e-09, 
    7.536277e-09, 8.041089e-09, 7.169219e-09, 7.654629e-09, 7.576224e-09, 
    8.058155e-09, 1.140321e-08, 1.070736e-08, 1.144544e-08, 1.134396e-08, 
    1.138943e-08, 1.195239e-08, 1.224362e-08, 1.287051e-08, 1.275502e-08, 
    1.229543e-08, 1.129855e-08, 1.16301e-08, 1.080802e-08, 1.08261e-08, 
    9.960975e-09, 1.034446e-08, 8.968475e-09, 9.344819e-09, 8.288354e-09, 
    8.545169e-09, 8.300276e-09, 8.373979e-09, 8.299319e-09, 8.678359e-09, 
    8.514405e-09, 8.853687e-09, 1.027181e-08, 9.838725e-09, 1.117175e-08, 
    1.203442e-08, 1.263387e-08, 1.307218e-08, 1.300955e-08, 1.289075e-08, 
    1.229278e-08, 1.174933e-08, 1.134712e-08, 1.108376e-08, 1.08287e-08, 
    1.008279e-08, 9.703871e-09, 8.89374e-09, 9.036126e-09, 8.795943e-09, 
    8.571042e-09, 8.203096e-09, 8.262836e-09, 8.103666e-09, 8.802256e-09, 
    8.333143e-09, 9.117974e-09, 8.898051e-09, 1.075988e-08, 1.153997e-08, 
    1.188358e-08, 1.219062e-08, 1.296154e-08, 1.242547e-08, 1.263482e-08, 
    1.214098e-08, 1.183457e-08, 1.198541e-08, 1.107662e-08, 1.142369e-08, 
    9.681748e-09, 1.040607e-08, 8.597049e-09, 9.006768e-09, 8.500957e-09, 
    8.756343e-09, 8.322176e-09, 8.712178e-09, 8.045035e-09, 7.904978e-09, 
    8.000484e-09, 7.638354e-09, 8.734185e-09, 8.300258e-09, 1.198965e-08, 
    1.196494e-08, 1.185037e-08, 1.236005e-08, 1.239175e-08, 1.287368e-08, 
    1.244423e-08, 1.226454e-08, 1.1817e-08, 1.155793e-08, 1.131555e-08, 
    1.079578e-08, 1.023626e-08, 9.49023e-09, 8.979774e-09, 8.649246e-09, 
    8.850837e-09, 8.672679e-09, 8.872009e-09, 8.966612e-09, 7.957227e-09, 
    8.512876e-09, 7.689664e-09, 7.73359e-09, 8.099902e-09, 7.728631e-09, 
    1.194762e-08, 1.209014e-08, 1.259451e-08, 1.219852e-08, 1.292697e-08, 
    1.251539e-08, 1.228309e-08, 1.141631e-08, 1.12321e-08, 1.106317e-08, 
    1.073508e-08, 1.032457e-08, 9.632588e-09, 9.059059e-09, 8.5581e-09, 
    8.594089e-09, 8.581404e-09, 8.47214e-09, 8.744689e-09, 8.428012e-09, 
    8.375697e-09, 8.512966e-09, 7.739486e-09, 7.954839e-09, 7.734526e-09, 
    7.874176e-09, 1.204368e-08, 1.180527e-08, 1.193366e-08, 1.169306e-08, 
    1.186217e-08, 1.112363e-08, 1.090894e-08, 9.944697e-09, 1.033253e-08, 
    9.720485e-09, 1.026911e-08, 1.017025e-08, 9.700892e-09, 1.02389e-08, 
    9.089963e-09, 9.857724e-09, 8.467914e-09, 9.195477e-09, 8.423798e-09, 
    8.560221e-09, 8.335256e-09, 8.13754e-09, 7.893865e-09, 7.458656e-09, 
    7.557791e-09, 7.204456e-09, 1.145631e-08, 1.115886e-08, 1.118487e-08, 
    1.087921e-08, 1.065713e-08, 1.018733e-08, 9.46599e-09, 9.732659e-09, 
    9.247335e-09, 9.152103e-09, 9.891135e-09, 9.432299e-09, 1.096302e-08, 
    1.070407e-08, 1.085773e-08, 1.143261e-08, 9.670663e-09, 1.054772e-08, 
    8.971505e-09, 9.41444e-09, 8.165509e-09, 8.770002e-09, 7.612778e-09, 
    7.159986e-09, 6.747237e-09, 6.288078e-09, 1.099899e-08, 1.119835e-08, 
    1.084328e-08, 1.03657e-08, 9.936758e-09, 9.386959e-09, 9.332032e-09, 
    9.232025e-09, 8.976739e-09, 8.766183e-09, 9.200533e-09, 8.713988e-09, 
    1.064458e-08, 9.597191e-09, 1.127437e-08, 1.074822e-08, 1.039344e-08, 
    1.054803e-08, 9.763499e-09, 9.585054e-09, 8.884726e-09, 9.241841e-09, 
    7.265783e-09, 8.096182e-09, 5.954995e-09, 6.505389e-09, 1.126862e-08, 
    1.099969e-08, 1.01004e-08, 1.052124e-08, 9.351101e-09, 9.078525e-09, 
    8.861373e-09, 8.589397e-09, 8.560439e-09, 8.402672e-09, 8.662349e-09, 
    8.412832e-09, 9.385813e-09, 8.94119e-09, 1.02004e-08, 9.882501e-09, 
    1.002783e-08, 1.018903e-08, 9.697608e-09, 9.193562e-09, 9.183075e-09, 
    9.02578e-09, 8.593226e-09, 9.346567e-09, 7.168642e-09, 8.459937e-09, 
    1.071185e-08, 1.021693e-08, 1.014773e-08, 1.033644e-08, 9.10558e-09, 
    9.538225e-09, 8.4065e-09, 8.701914e-09, 8.221869e-09, 8.457858e-09, 
    8.492998e-09, 8.804461e-09, 9.002615e-09, 9.518048e-09, 9.953355e-09, 
    1.030892e-08, 1.022542e-08, 9.837693e-09, 9.163392e-09, 8.557792e-09, 
    8.687807e-09, 8.257639e-09, 9.432534e-09, 8.925626e-09, 9.119058e-09, 
    8.621141e-09, 9.739806e-09, 8.780629e-09, 9.996953e-09, 9.8856e-09, 
    9.546965e-09, 8.891953e-09, 8.751778e-09, 8.603824e-09, 8.69491e-09, 
    9.146746e-09, 9.222435e-09, 9.555108e-09, 9.648476e-09, 9.90977e-09, 
    1.013e-08, 9.928626e-09, 9.720341e-09, 9.146579e-09, 8.651432e-09, 
    8.134743e-09, 8.011927e-09, 7.44443e-09, 7.903932e-09, 7.161838e-09, 
    7.788267e-09, 6.723984e-09, 8.727388e-09, 7.807575e-09, 9.531786e-09, 
    9.33356e-09, 8.982762e-09, 8.215534e-09, 8.623434e-09, 8.147886e-09, 
    9.225415e-09, 9.824479e-09, 9.984147e-09, 1.028702e-08, 9.977301e-09, 
    1.000223e-08, 9.711832e-09, 9.804467e-09, 9.127972e-09, 9.48689e-09, 
    8.493866e-09, 8.151577e-09, 7.240868e-09, 6.725934e-09, 6.22614e-09, 
    6.014789e-09, 5.951577e-09, 5.925302e-09,
  8.841753e-11, 8.066262e-11, 8.212644e-11, 7.618851e-11, 7.943886e-11, 
    7.561371e-11, 8.679988e-11, 8.036599e-11, 8.442803e-11, 8.769663e-11, 
    6.564503e-11, 7.593191e-11, 5.618732e-11, 6.185274e-11, 4.843884e-11, 
    5.703951e-11, 4.684304e-11, 4.867139e-11, 4.334439e-11, 4.481747e-11, 
    3.855546e-11, 4.267853e-11, 3.241818e-11, 3.950776e-11, 3.887589e-11, 
    4.282068e-11, 7.376499e-11, 6.686057e-11, 7.419118e-11, 7.316839e-11, 
    7.362608e-11, 7.937036e-11, 8.239683e-11, 8.90342e-11, 8.7799e-11, 
    8.293911e-11, 7.271219e-11, 7.606445e-11, 6.784522e-11, 6.802261e-11, 
    5.971313e-11, 6.335107e-11, 5.065151e-11, 5.402577e-11, 4.475515e-11, 
    4.695036e-11, 4.485621e-11, 4.548276e-11, 4.484809e-11, 4.810393e-11, 
    4.668537e-11, 4.963786e-11, 6.265624e-11, 5.856902e-11, 7.14433e-11, 
    8.021907e-11, 8.650927e-11, 9.120416e-11, 9.052849e-11, 8.925125e-11, 
    8.29113e-11, 7.728207e-11, 7.32001e-11, 7.056724e-11, 6.804814e-11, 
    6.086075e-11, 5.731588e-11, 4.999072e-11, 5.125234e-11, 4.913074e-11, 
    4.717365e-11, 4.403499e-11, 4.453915e-11, 4.32006e-11, 4.918609e-11, 
    4.513521e-11, 5.198263e-11, 5.002876e-11, 6.737367e-11, 7.514826e-11, 
    7.866068e-11, 8.184334e-11, 9.001164e-11, 8.430515e-11, 8.651942e-11, 
    8.132604e-11, 7.815651e-11, 7.971169e-11, 7.049633e-11, 7.397166e-11, 
    5.71112e-11, 6.394233e-11, 4.739849e-11, 5.099129e-11, 4.656971e-11, 
    4.878406e-11, 4.504204e-11, 4.839845e-11, 4.271138e-11, 4.155124e-11, 
    4.234105e-11, 3.937627e-11, 4.859045e-11, 4.485606e-11, 7.975549e-11, 
    7.950006e-11, 7.831891e-11, 8.3617e-11, 8.395026e-11, 8.906812e-11, 
    8.45028e-11, 8.261566e-11, 7.797605e-11, 7.533053e-11, 7.288283e-11, 
    6.772521e-11, 6.231715e-11, 5.535e-11, 5.075168e-11, 4.78509e-11, 
    4.961279e-11, 4.805452e-11, 4.979917e-11, 5.0635e-11, 4.198263e-11, 
    4.66722e-11, 3.979136e-11, 4.014804e-11, 4.316913e-11, 4.010772e-11, 
    7.932113e-11, 8.079726e-11, 8.609156e-11, 8.192571e-11, 8.964004e-11, 
    8.525397e-11, 8.280983e-11, 7.38971e-11, 7.204629e-11, 7.036276e-11, 
    6.713128e-11, 6.316058e-11, 5.665729e-11, 5.145659e-11, 4.706191e-11, 
    4.737287e-11, 4.726319e-11, 4.63222e-11, 4.868219e-11, 4.594414e-11, 
    4.549741e-11, 4.667299e-11, 4.019601e-11, 4.196288e-11, 4.015565e-11, 
    4.12977e-11, 8.031513e-11, 7.785562e-11, 7.917703e-11, 7.670665e-11, 
    7.844034e-11, 7.096381e-11, 6.883731e-11, 5.956034e-11, 6.323674e-11, 
    5.746976e-11, 6.263043e-11, 6.168932e-11, 5.72883e-11, 6.234236e-11, 
    5.173228e-11, 5.874633e-11, 4.628595e-11, 5.267754e-11, 4.590809e-11, 
    4.708021e-11, 4.515317e-11, 4.34842e-11, 4.14597e-11, 3.793577e-11, 
    3.87279e-11, 3.593381e-11, 7.430111e-11, 7.131483e-11, 7.157427e-11, 
    6.854456e-11, 6.637097e-11, 6.185153e-11, 5.512847e-11, 5.758261e-11, 
    5.314434e-11, 5.228823e-11, 5.905858e-11, 5.482108e-11, 6.937099e-11, 
    6.682844e-11, 6.833336e-11, 7.406168e-11, 5.700874e-11, 6.530886e-11, 
    5.067837e-11, 5.465838e-11, 4.371887e-11, 4.890353e-11, 3.916999e-11, 
    3.236421e-11, 2.996439e-11, 2.732572e-11, 6.972662e-11, 7.170891e-11, 
    6.819136e-11, 6.355474e-11, 5.948589e-11, 5.440837e-11, 5.390985e-11, 
    5.300637e-11, 5.072478e-11, 4.887012e-11, 5.272298e-11, 4.841423e-11, 
    6.624881e-11, 5.633123e-11, 7.246961e-11, 6.725966e-11, 6.382095e-11, 
    6.531187e-11, 5.786882e-11, 5.621959e-11, 4.991123e-11, 5.309481e-11, 
    3.64129e-11, 4.313803e-11, 2.543349e-11, 2.857033e-11, 7.241197e-11, 
    6.973359e-11, 6.102727e-11, 6.505266e-11, 5.408274e-11, 5.163019e-11, 
    4.970551e-11, 4.733229e-11, 4.70821e-11, 4.572755e-11, 4.796473e-11, 
    4.581435e-11, 5.439795e-11, 5.04099e-11, 6.197576e-11, 5.897784e-11, 
    6.034207e-11, 6.186771e-11, 5.725791e-11, 5.266033e-11, 5.256612e-11, 
    5.116029e-11, 4.73654e-11, 5.404162e-11, 3.24148e-11, 4.621753e-11, 
    6.690439e-11, 6.21331e-11, 6.147556e-11, 6.32742e-11, 5.187181e-11, 
    5.578955e-11, 4.576025e-11, 4.8309e-11, 4.419319e-11, 4.619971e-11, 
    4.65013e-11, 4.920543e-11, 5.09544e-11, 5.560461e-11, 5.964159e-11, 
    6.301079e-11, 6.221393e-11, 5.85594e-11, 5.238946e-11, 4.705925e-11, 
    4.818614e-11, 4.449521e-11, 5.482322e-11, 5.027226e-11, 5.199232e-11, 
    4.760711e-11, 5.764889e-11, 4.899656e-11, 6.005129e-11, 5.900681e-11, 
    5.586973e-11, 4.997495e-11, 4.874414e-11, 4.745712e-11, 4.824798e-11, 
    5.224022e-11, 5.292002e-11, 5.594446e-11, 5.680385e-11, 5.923299e-11, 
    6.130749e-11, 5.940964e-11, 5.746843e-11, 5.223872e-11, 4.786989e-11, 
    4.346075e-11, 4.243605e-11, 3.782262e-11, 4.154261e-11, 3.237503e-11, 
    4.05937e-11, 2.982995e-11, 4.853112e-11, 4.075152e-11, 5.573051e-11, 
    5.39237e-11, 5.077819e-11, 4.413978e-11, 4.762699e-11, 4.357095e-11, 
    5.294684e-11, 5.84362e-11, 5.993085e-11, 6.280151e-11, 5.986649e-11, 
    6.010098e-11, 5.73896e-11, 5.824979e-11, 5.207209e-11, 5.531946e-11, 
    4.650876e-11, 4.360192e-11, 3.621797e-11, 2.984122e-11, 2.697241e-11, 
    2.577176e-11, 2.541417e-11, 2.526575e-11,
  8.522608e-14, 7.269575e-14, 7.502895e-14, 6.566397e-14, 7.075725e-14, 
    6.477191e-14, 8.257871e-14, 7.222485e-14, 7.872833e-14, 8.404419e-14, 
    4.975649e-14, 6.526541e-14, 3.643887e-14, 4.429569e-14, 2.637755e-14, 
    3.759586e-14, 2.44193e-14, 2.666643e-14, 2.028254e-14, 2.199696e-14, 
    1.501375e-14, 1.952132e-14, 1.202253e-14, 1.602172e-14, 1.535057e-14, 
    1.968309e-14, 6.192114e-14, 5.153814e-14, 6.257583e-14, 6.100725e-14, 
    6.170808e-14, 7.064907e-14, 7.54616e-14, 8.623974e-14, 8.421181e-14, 
    7.633092e-14, 6.031047e-14, 6.54712e-14, 5.299198e-14, 5.325488e-14, 
    4.128389e-14, 4.643509e-14, 2.916089e-14, 3.354656e-14, 2.192362e-14, 
    2.454965e-14, 2.20426e-14, 2.278449e-14, 2.203304e-14, 2.596307e-14, 
    2.422815e-14, 2.787628e-14, 4.543995e-14, 3.969512e-14, 5.838192e-14, 
    7.199186e-14, 8.210491e-14, 8.982566e-14, 8.870597e-14, 8.65971e-14, 
    7.628629e-14, 6.736839e-14, 6.105575e-14, 5.705869e-14, 5.329274e-14, 
    4.289286e-14, 3.797303e-14, 2.832167e-14, 2.99297e-14, 2.72396e-14, 
    2.482149e-14, 2.108117e-14, 2.166992e-14, 2.011743e-14, 2.73089e-14, 
    2.237208e-14, 3.087139e-14, 2.836979e-14, 5.229456e-14, 6.405153e-14, 
    6.953042e-14, 7.457649e-14, 8.785136e-14, 7.852989e-14, 8.212144e-14, 
    7.375125e-14, 6.873805e-14, 7.118846e-14, 5.695189e-14, 6.223841e-14, 
    3.76936e-14, 4.728594e-14, 2.509607e-14, 2.959501e-14, 2.40882e-14, 
    2.68067e-14, 2.226189e-14, 2.632747e-14, 1.955867e-14, 1.825283e-14, 
    1.913886e-14, 1.588132e-14, 2.656579e-14, 2.204242e-14, 7.125774e-14, 
    7.085393e-14, 6.899306e-14, 7.742053e-14, 7.795736e-14, 8.629557e-14, 
    7.884913e-14, 7.581217e-14, 6.845489e-14, 6.433343e-14, 6.05709e-14, 
    5.281429e-14, 4.49562e-14, 3.531115e-14, 2.928869e-14, 2.565114e-14, 
    2.784472e-14, 2.590207e-14, 2.807965e-14, 2.913984e-14, 1.873519e-14, 
    2.421221e-14, 1.632591e-14, 1.671101e-14, 2.008134e-14, 1.666733e-14, 
    7.057136e-14, 7.29097e-14, 8.14249e-14, 7.470809e-14, 8.723796e-14, 
    8.006483e-14, 7.612348e-14, 6.212392e-14, 5.929664e-14, 5.675083e-14, 
    5.19369e-14, 4.616176e-14, 3.707579e-14, 3.019228e-14, 2.468535e-14, 
    2.506474e-14, 2.493073e-14, 2.378951e-14, 2.667987e-14, 2.333533e-14, 
    2.280193e-14, 2.421316e-14, 1.676302e-14, 1.871303e-14, 1.671926e-14, 
    1.797115e-14, 7.214417e-14, 6.826608e-14, 7.034397e-14, 6.647035e-14, 
    6.91839e-14, 5.765683e-14, 5.446618e-14, 4.107083e-14, 4.627099e-14, 
    3.818346e-14, 4.540308e-14, 4.406384e-14, 3.793535e-14, 4.499212e-14, 
    3.054769e-14, 3.994031e-14, 2.374585e-14, 3.177464e-14, 2.329216e-14, 
    2.470763e-14, 2.239334e-14, 2.044348e-14, 1.815098e-14, 1.436922e-14, 
    1.519472e-14, 1.23516e-14, 6.274493e-14, 5.818744e-14, 5.858031e-14, 
    5.403019e-14, 5.081876e-14, 4.429398e-14, 3.501432e-14, 3.833797e-14, 
    3.238527e-14, 3.126776e-14, 4.037305e-14, 3.460353e-14, 5.526302e-14, 
    5.149085e-14, 5.371616e-14, 6.237674e-14, 3.755393e-14, 4.926636e-14, 
    2.919515e-14, 3.438661e-14, 2.071447e-14, 2.695567e-14, 1.566182e-14, 
    1.195312e-14, 9.047565e-15, 6.281994e-15, 5.579549e-14, 5.878444e-14, 
    5.350527e-14, 4.672775e-14, 4.09671e-14, 3.405397e-14, 3.339323e-14, 
    3.220447e-14, 2.925435e-14, 2.691399e-14, 3.183395e-14, 2.634703e-14, 
    5.063962e-14, 3.66336e-14, 5.99407e-14, 5.212627e-14, 4.711096e-14, 
    4.927076e-14, 3.873053e-14, 3.648251e-14, 2.822116e-14, 3.232033e-14, 
    1.282519e-14, 2.00457e-14, 4.59418e-15, 7.528406e-15, 5.985291e-14, 
    5.580593e-14, 4.312759e-14, 4.889363e-14, 3.3622e-14, 3.041595e-14, 
    2.796152e-14, 2.501513e-14, 2.470993e-14, 2.307628e-14, 2.579132e-14, 
    2.317999e-14, 3.404013e-14, 2.885327e-14, 4.447044e-14, 4.026104e-14, 
    4.216381e-14, 4.431695e-14, 3.789385e-14, 3.17522e-14, 3.162935e-14, 
    2.981156e-14, 2.50556e-14, 3.356755e-14, 1.201818e-14, 2.366352e-14, 
    5.160264e-14, 4.469416e-14, 4.376102e-14, 4.632473e-14, 3.072799e-14, 
    3.590201e-14, 2.311533e-14, 2.621664e-14, 2.12654e-14, 2.364209e-14, 
    2.400554e-14, 2.733313e-14, 2.954779e-14, 3.56531e-14, 4.118409e-14, 
    4.59471e-14, 4.480919e-14, 3.968183e-14, 3.139935e-14, 2.468211e-14, 
    2.606464e-14, 2.161841e-14, 3.460639e-14, 2.867842e-14, 3.088394e-14, 
    2.53516e-14, 3.842879e-14, 2.707183e-14, 4.175641e-14, 4.030123e-14, 
    3.601006e-14, 2.830173e-14, 2.675699e-14, 2.516781e-14, 2.614112e-14, 
    3.12054e-14, 3.209145e-14, 3.611084e-14, 3.727499e-14, 4.061525e-14, 
    4.352327e-14, 4.086094e-14, 3.818164e-14, 3.120345e-14, 2.567451e-14, 
    2.041647e-14, 1.924629e-14, 1.425253e-14, 1.824323e-14, 1.196702e-14, 
    1.719611e-14, 8.895531e-15, 2.649207e-14, 1.736894e-14, 3.58225e-14, 
    3.341155e-14, 2.932253e-14, 2.120315e-14, 2.537599e-14, 2.054353e-14, 
    3.212655e-14, 3.951169e-14, 4.158797e-14, 4.564758e-14, 4.149803e-14, 
    4.182596e-14, 3.807381e-14, 3.925461e-14, 3.098728e-14, 3.52702e-14, 
    2.401455e-14, 2.057929e-14, 1.263177e-14, 8.908233e-15, 5.947605e-15, 
    4.877095e-15, 4.578274e-15, 4.456975e-15,
  2.880587e-19, 2.462414e-19, 2.540361e-19, 2.227253e-19, 2.397623e-19, 
    2.197393e-19, 2.792324e-19, 2.446677e-19, 2.663871e-19, 2.841189e-19, 
    1.693738e-19, 2.213912e-19, 1.245086e-19, 1.510022e-19, 9.045994e-20, 
    1.28415e-19, 8.381285e-20, 9.143987e-20, 6.974473e-20, 7.557966e-20, 
    5.176569e-20, 6.715172e-20, 4.156026e-20, 5.521132e-20, 5.291743e-20, 
    6.770289e-20, 2.101924e-19, 1.753609e-19, 2.123855e-19, 2.071305e-19, 
    2.094787e-19, 2.394006e-19, 2.554811e-19, 2.914371e-19, 2.846777e-19, 
    2.58384e-19, 2.047955e-19, 2.220801e-19, 1.802441e-19, 1.811269e-19, 
    1.408553e-19, 1.582035e-19, 9.989536e-20, 1.14736e-19, 7.533016e-20, 
    8.425554e-20, 7.573488e-20, 7.825774e-20, 7.570235e-20, 8.905363e-20, 
    8.31636e-20, 9.554233e-20, 1.548545e-19, 1.354982e-19, 1.983305e-19, 
    2.438891e-19, 2.776523e-19, 3.033833e-19, 2.99654e-19, 2.92628e-19, 
    2.58235e-19, 2.284288e-19, 2.07293e-19, 1.938928e-19, 1.812541e-19, 
    1.462773e-19, 1.29688e-19, 9.705189e-20, 1.024992e-19, 9.338377e-20, 
    8.517865e-20, 7.246365e-20, 7.44671e-20, 6.918239e-20, 9.361874e-20, 
    7.685546e-20, 1.056872e-19, 9.721498e-20, 1.779019e-19, 2.173275e-19, 
    2.356604e-19, 2.525249e-19, 2.968071e-19, 2.657248e-19, 2.777074e-19, 
    2.497681e-19, 2.330104e-19, 2.412038e-19, 1.935345e-19, 2.112553e-19, 
    1.287449e-19, 1.610662e-19, 8.611092e-20, 1.013658e-19, 8.268822e-20, 
    9.191567e-20, 7.648073e-20, 9.029002e-20, 6.727896e-20, 6.282754e-20, 
    6.584836e-20, 5.473155e-20, 9.109851e-20, 7.573427e-20, 2.414354e-19, 
    2.400855e-19, 2.338634e-19, 2.620219e-19, 2.638139e-19, 2.916231e-19, 
    2.667903e-19, 2.566518e-19, 2.320634e-19, 2.182713e-19, 2.056683e-19, 
    1.796474e-19, 1.53226e-19, 1.206993e-19, 1.003283e-19, 8.799508e-20, 
    9.543532e-20, 8.884664e-20, 9.623165e-20, 9.982408e-20, 6.447236e-20, 
    8.310947e-20, 5.625054e-20, 5.756581e-20, 6.905949e-20, 5.741664e-20, 
    2.391408e-19, 2.469563e-19, 2.753842e-19, 2.529644e-19, 2.947634e-19, 
    2.70847e-19, 2.576914e-19, 2.108717e-19, 2.013973e-19, 1.928601e-19, 
    1.767005e-19, 1.572838e-19, 1.266593e-19, 1.033883e-19, 8.471636e-20, 
    8.600457e-20, 8.554958e-20, 8.167347e-20, 9.148547e-20, 8.013012e-20, 
    7.831701e-20, 8.31127e-20, 5.77434e-20, 6.439678e-20, 5.759397e-20, 
    6.186674e-20, 2.443981e-19, 2.314318e-19, 2.383806e-19, 2.25424e-19, 
    2.345016e-19, 1.95899e-19, 1.851936e-19, 1.401371e-19, 1.576514e-19, 
    1.303982e-19, 1.547304e-19, 1.502215e-19, 1.295609e-19, 1.53347e-19, 
    1.045915e-19, 1.363252e-19, 8.152513e-20, 1.087437e-19, 7.99834e-20, 
    8.479204e-20, 7.692776e-20, 7.029277e-20, 6.248015e-20, 4.956077e-20, 
    5.238455e-20, 4.264936e-20, 2.129519e-19, 1.976784e-19, 1.989957e-19, 
    1.8373e-19, 1.729439e-19, 1.509964e-19, 1.196963e-19, 1.309196e-19, 
    1.108093e-19, 1.070286e-19, 1.377845e-19, 1.183082e-19, 1.878681e-19, 
    1.75202e-19, 1.826758e-19, 2.117186e-19, 1.282734e-19, 1.677262e-19, 
    1.000114e-19, 1.175752e-19, 7.121539e-20, 9.242091e-20, 5.39814e-20, 
    4.132195e-20, 3.132731e-20, 2.177434e-20, 1.896549e-19, 1.996801e-19, 
    1.819677e-19, 1.591883e-19, 1.397874e-19, 1.164511e-19, 1.142177e-19, 
    1.101978e-19, 1.002119e-19, 9.227955e-20, 1.089444e-19, 9.03564e-20, 
    1.723419e-19, 1.251662e-19, 2.035562e-19, 1.773366e-19, 1.604775e-19, 
    1.677409e-19, 1.322442e-19, 1.24656e-19, 9.671127e-20, 1.105897e-19, 
    4.427294e-20, 6.893811e-20, 1.591863e-20, 2.608519e-20, 2.032619e-19, 
    1.896899e-19, 1.470681e-19, 1.66473e-19, 1.14991e-19, 1.041455e-19, 
    9.583123e-20, 8.583613e-20, 8.479984e-20, 7.924964e-20, 8.847084e-20, 
    7.960216e-20, 1.164043e-19, 9.88532e-20, 1.515906e-19, 1.374068e-19, 
    1.438209e-19, 1.510738e-19, 1.294208e-19, 1.086678e-19, 1.082522e-19, 
    1.020992e-19, 8.597353e-20, 1.14807e-19, 4.154534e-20, 8.124538e-20, 
    1.755776e-19, 1.523438e-19, 1.492016e-19, 1.578322e-19, 1.052018e-19, 
    1.226954e-19, 7.938237e-20, 8.991402e-20, 7.309064e-20, 8.117257e-20, 
    8.240741e-20, 9.370089e-20, 1.012059e-19, 1.218545e-19, 1.405189e-19, 
    1.565614e-19, 1.527311e-19, 1.354534e-19, 1.074739e-19, 8.470537e-20, 
    8.939828e-20, 7.429186e-20, 1.183178e-19, 9.826078e-20, 1.057297e-19, 
    8.69784e-20, 1.312261e-19, 9.281484e-20, 1.42448e-19, 1.375423e-19, 
    1.230603e-19, 9.69843e-20, 9.174705e-20, 8.635446e-20, 8.965779e-20, 
    1.068176e-19, 1.098155e-19, 1.234007e-19, 1.273318e-19, 1.386011e-19, 
    1.484009e-19, 1.394295e-19, 1.303921e-19, 1.06811e-19, 8.807439e-20, 
    7.020077e-20, 6.621452e-20, 4.916141e-20, 6.279478e-20, 4.136968e-20, 
    5.9222e-20, 3.080325e-20, 9.084845e-20, 5.98119e-20, 1.224268e-19, 
    1.142796e-19, 1.004429e-19, 7.287879e-20, 8.706117e-20, 7.063342e-20, 
    1.099342e-19, 1.348795e-19, 1.418802e-19, 1.555533e-19, 1.415771e-19, 
    1.426823e-19, 1.300282e-19, 1.340123e-19, 1.060795e-19, 1.205609e-19, 
    8.243801e-20, 7.075516e-20, 4.360996e-20, 3.084704e-20, 2.061602e-20, 
    1.690186e-20, 1.586333e-20, 1.544152e-20,
  2.114393e-25, 1.808953e-25, 1.865904e-25, 1.637085e-25, 1.761608e-25, 
    1.615256e-25, 2.049942e-25, 1.797454e-25, 1.956128e-25, 2.085625e-25, 
    1.246823e-25, 1.627333e-25, 9.181547e-26, 1.112302e-25, 6.682709e-26, 
    9.467938e-26, 6.194306e-26, 6.754692e-26, 5.159872e-26, 5.589052e-26, 
    3.835989e-26, 4.96908e-26, 3.0843e-26, 4.089902e-26, 3.920874e-26, 
    5.009638e-26, 1.545454e-25, 1.290646e-25, 1.56149e-25, 1.523063e-25, 
    1.540234e-25, 1.758965e-25, 1.87646e-25, 2.13906e-25, 2.089705e-25, 
    1.897667e-25, 1.505987e-25, 1.632368e-25, 1.326383e-25, 1.332843e-25, 
    1.037968e-25, 1.165041e-25, 7.375642e-26, 8.464818e-26, 5.570705e-26, 
    6.22684e-26, 5.600467e-26, 5.785968e-26, 5.598075e-26, 6.579396e-26, 
    6.14659e-26, 7.056005e-26, 1.140516e-25, 9.98712e-26, 1.458704e-25, 
    1.791765e-25, 2.038403e-25, 2.226275e-25, 2.19905e-25, 2.147755e-25, 
    1.896579e-25, 1.678777e-25, 1.524252e-25, 1.426243e-25, 1.333773e-25, 
    1.077692e-25, 9.561262e-26, 7.166859e-26, 7.566802e-26, 6.897474e-26, 
    6.294677e-26, 5.359885e-26, 5.507235e-26, 5.1185e-26, 6.914733e-26, 
    5.682865e-26, 7.800813e-26, 7.178835e-26, 1.309242e-25, 1.597623e-25, 
    1.731631e-25, 1.854863e-25, 2.178266e-25, 1.95129e-25, 2.038805e-25, 
    1.834721e-25, 1.712264e-25, 1.772142e-25, 1.423622e-25, 1.553225e-25, 
    9.492124e-26, 1.186002e-25, 6.363184e-26, 7.483594e-26, 6.111652e-26, 
    6.789642e-26, 5.655312e-26, 6.670226e-26, 4.978443e-26, 4.650808e-26, 
    4.873162e-26, 4.054552e-26, 6.729617e-26, 5.600422e-26, 1.773835e-25, 
    1.76397e-25, 1.718498e-25, 1.924242e-25, 1.937332e-25, 2.140419e-25, 
    1.959072e-25, 1.885013e-25, 1.705342e-25, 1.604523e-25, 1.51237e-25, 
    1.322016e-25, 1.12859e-25, 8.902225e-26, 7.407427e-26, 6.501625e-26, 
    7.048146e-26, 6.564189e-26, 7.106626e-26, 7.370409e-26, 4.771887e-26, 
    6.142612e-26, 4.166463e-26, 4.263349e-26, 5.109457e-26, 4.252362e-26, 
    1.757067e-25, 1.814177e-25, 2.021839e-25, 1.858074e-25, 2.163345e-25, 
    1.988702e-25, 1.892607e-25, 1.550421e-25, 1.481135e-25, 1.418688e-25, 
    1.30045e-25, 1.158306e-25, 9.339226e-26, 7.632068e-26, 6.260705e-26, 
    6.355369e-26, 6.321936e-26, 6.037067e-26, 6.758042e-26, 5.923619e-26, 
    5.790327e-26, 6.142849e-26, 4.27643e-26, 4.766324e-26, 4.265424e-26, 
    4.580073e-26, 1.795484e-25, 1.700727e-25, 1.751511e-25, 1.656813e-25, 
    1.723162e-25, 1.440918e-25, 1.3626e-25, 1.032705e-25, 1.160998e-25, 
    9.613319e-26, 1.139607e-25, 1.106583e-25, 9.551939e-26, 1.129475e-25, 
    7.720389e-26, 1.004772e-25, 6.026163e-26, 8.025134e-26, 5.912834e-26, 
    6.266267e-26, 5.688181e-26, 5.200191e-26, 4.625234e-26, 3.67345e-26, 
    3.881601e-26, 3.163655e-26, 1.565631e-25, 1.453934e-25, 1.463569e-25, 
    1.351891e-25, 1.272955e-25, 1.112259e-25, 8.828674e-26, 9.651539e-26, 
    8.176709e-26, 7.899266e-26, 1.015466e-25, 8.726867e-26, 1.382168e-25, 
    1.289483e-25, 1.344176e-25, 1.556613e-25, 9.457562e-26, 1.234762e-25, 
    7.384162e-26, 8.6731e-26, 5.268064e-26, 6.826753e-26, 3.999279e-26, 
    3.066704e-26, 2.3281e-26, 1.620576e-26, 1.39524e-25, 1.468575e-25, 
    1.338995e-25, 1.172252e-25, 1.030143e-25, 8.590637e-26, 8.426789e-26, 
    8.131836e-26, 7.398885e-26, 6.81637e-26, 8.039858e-26, 6.675102e-26, 
    1.268549e-25, 9.229763e-26, 1.496924e-25, 1.305105e-25, 1.181692e-25, 
    1.23487e-25, 9.748632e-26, 9.192353e-26, 7.141846e-26, 8.160593e-26, 
    3.283457e-26, 5.100526e-26, 1.185807e-26, 1.940088e-26, 1.494772e-25, 
    1.395496e-25, 1.083484e-25, 1.225588e-25, 8.483525e-26, 7.687654e-26, 
    7.077221e-26, 6.342991e-26, 6.26684e-26, 5.858892e-26, 6.536579e-26, 
    5.884807e-26, 8.587206e-26, 7.299125e-26, 1.116612e-25, 1.012698e-25, 
    1.059696e-25, 1.112826e-25, 9.541669e-26, 8.019561e-26, 7.98906e-26, 
    7.537435e-26, 6.353088e-26, 8.470022e-26, 3.083199e-26, 6.0056e-26, 
    1.292231e-25, 1.122128e-25, 1.099113e-25, 1.162322e-25, 7.765186e-26, 
    9.048596e-26, 5.86865e-26, 6.642604e-26, 5.406001e-26, 6.000248e-26, 
    6.091012e-26, 6.920766e-26, 7.471854e-26, 8.98694e-26, 1.035503e-25, 
    1.153016e-25, 1.124965e-25, 9.983835e-26, 7.931945e-26, 6.259898e-26, 
    6.604716e-26, 5.494348e-26, 8.727575e-26, 7.255627e-26, 7.803929e-26, 
    6.426925e-26, 9.674003e-26, 6.855688e-26, 1.049637e-25, 1.013692e-25, 
    9.075356e-26, 7.161896e-26, 6.777256e-26, 6.381079e-26, 6.623781e-26, 
    7.883779e-26, 8.103782e-26, 9.100317e-26, 9.388529e-26, 1.021451e-25, 
    1.093248e-25, 1.027521e-25, 9.612869e-26, 7.883295e-26, 6.507452e-26, 
    5.193423e-26, 4.90011e-26, 3.644006e-26, 4.648397e-26, 3.070229e-26, 
    4.385329e-26, 2.289332e-26, 6.711248e-26, 4.428771e-26, 9.028901e-26, 
    8.431331e-26, 7.415842e-26, 5.390419e-26, 6.433007e-26, 5.225252e-26, 
    8.112494e-26, 9.941777e-26, 1.045478e-25, 1.145634e-25, 1.043257e-25, 
    1.051354e-25, 9.586194e-26, 9.87822e-26, 7.8296e-26, 8.892078e-26, 
    6.093261e-26, 5.234208e-26, 3.23454e-26, 2.292571e-26, 1.534649e-26, 
    1.25888e-26, 1.181696e-26, 1.150337e-26,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_SAT =
  0.0111753, 0.01118969, 0.01118689, 0.01119848, 0.01119205, 0.01119964, 
    0.01117821, 0.01119026, 0.01118257, 0.01117658, 0.01122093, 0.01119899, 
    0.01124355, 0.01122964, 0.01126454, 0.0112414, 0.01126919, 0.01126385, 
    0.01127986, 0.01127528, 0.01129573, 0.01128197, 0.01130628, 0.01129244, 
    0.01129462, 0.01128152, 0.0112034, 0.01121821, 0.01120252, 0.01120464, 
    0.01120369, 0.01119218, 0.01118639, 0.01117419, 0.0111764, 0.01118536, 
    0.01120559, 0.01119872, 0.01121598, 0.01121559, 0.01123477, 0.01122613, 
    0.01125827, 0.01124913, 0.01127547, 0.01126886, 0.01127516, 0.01127325, 
    0.01127519, 0.01126549, 0.01126965, 0.0112611, 0.01122775, 0.01123757, 
    0.01120824, 0.01119056, 0.01117874, 0.01117035, 0.01117154, 0.01117381, 
    0.01118541, 0.01119628, 0.01120456, 0.01121009, 0.01121554, 0.01123203, 
    0.0112407, 0.01126012, 0.0112566, 0.01126255, 0.0112682, 0.0112777, 
    0.01127614, 0.01128032, 0.01126238, 0.01127431, 0.0112546, 0.01126, 
    0.01121708, 0.01120057, 0.01119359, 0.01118743, 0.01117245, 0.0111828, 
    0.01117873, 0.0111884, 0.01119455, 0.01119151, 0.01121025, 0.01120297, 
    0.01124121, 0.01122477, 0.01126754, 0.01125732, 0.01126999, 0.01126353, 
    0.0112746, 0.01126463, 0.01128187, 0.01128562, 0.01128306, 0.01129288, 
    0.01126408, 0.01127517, 0.01119143, 0.01119193, 0.01119423, 0.01118409, 
    0.01118346, 0.01117413, 0.01118243, 0.01118596, 0.01119491, 0.0112002, 
    0.01120522, 0.01121625, 0.01122855, 0.01124569, 0.01125799, 0.01126622, 
    0.01126117, 0.01126563, 0.01126064, 0.0112583, 0.01128422, 0.01126969, 
    0.01129147, 0.01129026, 0.01128042, 0.0112904, 0.01119227, 0.01118942, 
    0.0111795, 0.01118726, 0.01117311, 0.01118104, 0.0111856, 0.01120314, 
    0.01120697, 0.01121054, 0.01121756, 0.01122657, 0.01124235, 0.01125605, 
    0.01126853, 0.01126761, 0.01126793, 0.01127073, 0.01126382, 0.01127186, 
    0.01127321, 0.01126968, 0.0112901, 0.01128428, 0.01129024, 0.01128644, 
    0.01119034, 0.01119515, 0.01119255, 0.01119743, 0.011194, 0.01120927, 
    0.01121384, 0.01123515, 0.0112264, 0.01124031, 0.01122781, 0.01123003, 
    0.01124078, 0.01122848, 0.0112553, 0.01123715, 0.01127083, 0.01125275, 
    0.01127197, 0.01126847, 0.01127425, 0.01127942, 0.01128592, 0.01129789, 
    0.01129512, 0.01130511, 0.0112023, 0.01120852, 0.01120796, 0.01121446, 
    0.01121926, 0.01122964, 0.01124626, 0.01124001, 0.01125147, 0.01125378, 
    0.01123636, 0.01124706, 0.01121267, 0.01121825, 0.01121492, 0.01120279, 
    0.01124147, 0.01122166, 0.01125819, 0.01124748, 0.01127869, 0.0112632, 
    0.01129359, 0.01130656, 0.01131869, 0.01133288, 0.0112119, 0.01120767, 
    0.01121522, 0.01122567, 0.01123532, 0.01124813, 0.01124944, 0.01125184, 
    0.01125806, 0.01126328, 0.01125261, 0.01126459, 0.01121957, 0.01124318, 
    0.01120609, 0.0112173, 0.01122505, 0.01122164, 0.01123929, 0.01124345, 
    0.01126034, 0.0112516, 0.01130337, 0.01128053, 0.01134363, 0.01132608, 
    0.0112062, 0.01121188, 0.01123161, 0.01122223, 0.01124898, 0.01125557, 
    0.01126091, 0.01126774, 0.01126847, 0.01127251, 0.01126589, 0.01127225, 
    0.01124816, 0.01125894, 0.01122934, 0.01123656, 0.01123324, 0.0112296, 
    0.01124082, 0.01125279, 0.01125302, 0.01125686, 0.0112677, 0.01124909, 
    0.01130635, 0.01127109, 0.01121806, 0.01122899, 0.01123053, 0.0112263, 
    0.01125491, 0.01124456, 0.01127241, 0.01126489, 0.0112772, 0.01127109, 
    0.01127019, 0.01126232, 0.01125742, 0.01124503, 0.01123494, 0.01122691, 
    0.01122878, 0.01123759, 0.01125351, 0.01126854, 0.01126526, 0.01127627, 
    0.01124705, 0.01125933, 0.01125459, 0.01126693, 0.01123985, 0.01126297, 
    0.01123394, 0.01123648, 0.01124435, 0.01126017, 0.01126364, 0.01126738, 
    0.01126507, 0.01125391, 0.01125208, 0.01124415, 0.01124198, 0.01123593, 
    0.01123092, 0.0112355, 0.01124031, 0.01125391, 0.01126617, 0.0112795, 
    0.01128275, 0.01129832, 0.01128567, 0.01130655, 0.01128884, 0.01131943, 
    0.01126428, 0.01128828, 0.0112447, 0.0112494, 0.01125793, 0.01127739, 
    0.01126687, 0.01127916, 0.011252, 0.0112379, 0.01123423, 0.01122741, 
    0.01123439, 0.01123382, 0.01124049, 0.01123835, 0.01125436, 0.01124576, 
    0.01127017, 0.01127906, 0.01130407, 0.01131935, 0.01133483, 0.01134166, 
    0.01134373, 0.0113446,
  3.669827e-05, 3.678982e-05, 3.6772e-05, 3.684585e-05, 3.680484e-05, 
    3.685322e-05, 3.671678e-05, 3.679351e-05, 3.67445e-05, 3.670644e-05, 
    3.698913e-05, 3.684912e-05, 3.71337e-05, 3.704471e-05, 3.726805e-05, 
    3.711994e-05, 3.729786e-05, 3.726364e-05, 3.736626e-05, 3.733687e-05, 
    3.746823e-05, 3.737981e-05, 3.7536e-05, 3.744705e-05, 3.746103e-05, 
    3.737692e-05, 3.687719e-05, 3.697176e-05, 3.687161e-05, 3.68851e-05, 
    3.687902e-05, 3.680574e-05, 3.676887e-05, 3.669118e-05, 3.670526e-05, 
    3.676227e-05, 3.689116e-05, 3.684734e-05, 3.695746e-05, 3.695497e-05, 
    3.707746e-05, 3.702226e-05, 3.722785e-05, 3.716937e-05, 3.733809e-05, 
    3.729572e-05, 3.733613e-05, 3.732386e-05, 3.733629e-05, 3.727413e-05, 
    3.730078e-05, 3.724601e-05, 3.703262e-05, 3.70954e-05, 3.690809e-05, 
    3.679543e-05, 3.672018e-05, 3.666683e-05, 3.667437e-05, 3.668878e-05, 
    3.676261e-05, 3.683184e-05, 3.688459e-05, 3.691988e-05, 3.695461e-05, 
    3.706e-05, 3.711543e-05, 3.723973e-05, 3.721719e-05, 3.725529e-05, 
    3.72915e-05, 3.735241e-05, 3.734237e-05, 3.736922e-05, 3.725419e-05, 
    3.733071e-05, 3.720437e-05, 3.723896e-05, 3.696452e-05, 3.685915e-05, 
    3.681471e-05, 3.677544e-05, 3.668018e-05, 3.674601e-05, 3.672007e-05, 
    3.678165e-05, 3.682082e-05, 3.680143e-05, 3.692084e-05, 3.687446e-05, 
    3.711872e-05, 3.70136e-05, 3.728728e-05, 3.72218e-05, 3.730294e-05, 
    3.726153e-05, 3.733251e-05, 3.726863e-05, 3.737917e-05, 3.740328e-05, 
    3.738682e-05, 3.744986e-05, 3.72651e-05, 3.733617e-05, 3.680091e-05, 
    3.680408e-05, 3.681877e-05, 3.675418e-05, 3.67502e-05, 3.669082e-05, 
    3.674362e-05, 3.676613e-05, 3.682305e-05, 3.68568e-05, 3.688882e-05, 
    3.695918e-05, 3.703776e-05, 3.714738e-05, 3.722605e-05, 3.727878e-05, 
    3.724642e-05, 3.7275e-05, 3.724307e-05, 3.722808e-05, 3.739428e-05, 
    3.730105e-05, 3.744079e-05, 3.743305e-05, 3.736988e-05, 3.743393e-05, 
    3.680629e-05, 3.678809e-05, 3.672501e-05, 3.677438e-05, 3.668434e-05, 
    3.673481e-05, 3.676385e-05, 3.687553e-05, 3.689994e-05, 3.69227e-05, 
    3.696753e-05, 3.702509e-05, 3.712598e-05, 3.721365e-05, 3.729359e-05, 
    3.728773e-05, 3.728979e-05, 3.730768e-05, 3.726342e-05, 3.731495e-05, 
    3.732363e-05, 3.730098e-05, 3.743202e-05, 3.73946e-05, 3.743289e-05, 
    3.740852e-05, 3.679399e-05, 3.68246e-05, 3.680807e-05, 3.683917e-05, 
    3.68173e-05, 3.691463e-05, 3.694379e-05, 3.707995e-05, 3.702398e-05, 
    3.71129e-05, 3.703298e-05, 3.704717e-05, 3.7116e-05, 3.703727e-05, 
    3.720891e-05, 3.709274e-05, 3.730838e-05, 3.71926e-05, 3.731564e-05, 
    3.729324e-05, 3.733027e-05, 3.736347e-05, 3.740513e-05, 3.748206e-05, 
    3.746423e-05, 3.752843e-05, 3.687015e-05, 3.690984e-05, 3.690626e-05, 
    3.694771e-05, 3.697837e-05, 3.704467e-05, 3.715099e-05, 3.7111e-05, 
    3.718434e-05, 3.71991e-05, 3.708761e-05, 3.715614e-05, 3.693632e-05, 
    3.697197e-05, 3.695068e-05, 3.687333e-05, 3.712034e-05, 3.699373e-05, 
    3.722737e-05, 3.715879e-05, 3.735875e-05, 3.725947e-05, 3.745444e-05, 
    3.753783e-05, 3.76158e-05, 3.770728e-05, 3.693139e-05, 3.690444e-05, 
    3.695261e-05, 3.701936e-05, 3.708099e-05, 3.716298e-05, 3.717133e-05, 
    3.718673e-05, 3.722649e-05, 3.725996e-05, 3.719168e-05, 3.726834e-05, 
    3.698041e-05, 3.713128e-05, 3.689433e-05, 3.696588e-05, 3.701538e-05, 
    3.699358e-05, 3.710641e-05, 3.7133e-05, 3.724114e-05, 3.718518e-05, 
    3.751734e-05, 3.737061e-05, 3.777654e-05, 3.766343e-05, 3.689505e-05, 
    3.693126e-05, 3.705726e-05, 3.699732e-05, 3.716841e-05, 3.721057e-05, 
    3.724475e-05, 3.728856e-05, 3.729322e-05, 3.731915e-05, 3.727666e-05, 
    3.731744e-05, 3.716316e-05, 3.723213e-05, 3.704277e-05, 3.708893e-05, 
    3.706766e-05, 3.70444e-05, 3.711619e-05, 3.719278e-05, 3.719428e-05, 
    3.721887e-05, 3.728837e-05, 3.71691e-05, 3.753651e-05, 3.73101e-05, 
    3.697073e-05, 3.704058e-05, 3.705038e-05, 3.702336e-05, 3.720635e-05, 
    3.714007e-05, 3.73185e-05, 3.727028e-05, 3.734923e-05, 3.731002e-05, 
    3.730426e-05, 3.725383e-05, 3.722246e-05, 3.714314e-05, 3.707857e-05, 
    3.702726e-05, 3.703919e-05, 3.709553e-05, 3.719743e-05, 3.729371e-05, 
    3.727265e-05, 3.734323e-05, 3.715602e-05, 3.723465e-05, 3.720431e-05, 
    3.728336e-05, 3.710997e-05, 3.725807e-05, 3.707215e-05, 3.708843e-05, 
    3.713876e-05, 3.724008e-05, 3.726227e-05, 3.728621e-05, 3.727141e-05, 
    3.72e-05, 3.718823e-05, 3.71375e-05, 3.712357e-05, 3.708487e-05, 
    3.705289e-05, 3.708215e-05, 3.71129e-05, 3.719997e-05, 3.72785e-05, 
    3.736397e-05, 3.738481e-05, 3.748485e-05, 3.740362e-05, 3.75378e-05, 
    3.742403e-05, 3.762068e-05, 3.726643e-05, 3.74204e-05, 3.7141e-05, 
    3.717108e-05, 3.722569e-05, 3.735047e-05, 3.728299e-05, 3.736183e-05, 
    3.718775e-05, 3.709755e-05, 3.707403e-05, 3.703041e-05, 3.707502e-05, 
    3.707139e-05, 3.711407e-05, 3.710035e-05, 3.720286e-05, 3.714778e-05, 
    3.730415e-05, 3.736117e-05, 3.752176e-05, 3.762008e-05, 3.771978e-05, 
    3.776381e-05, 3.77772e-05, 3.77828e-05,
  8.81479e-10, 8.842221e-10, 8.836878e-10, 8.859022e-10, 8.846723e-10, 
    8.861233e-10, 8.820333e-10, 8.843326e-10, 8.828638e-10, 8.817234e-10, 
    8.902034e-10, 8.860004e-10, 8.946326e-10, 8.918731e-10, 8.988095e-10, 
    8.942049e-10, 8.997371e-10, 8.986721e-10, 9.018662e-10, 9.00951e-10, 
    9.050443e-10, 9.022885e-10, 9.071581e-10, 9.043838e-10, 9.048196e-10, 
    9.021983e-10, 8.868423e-10, 8.896816e-10, 8.866751e-10, 8.870797e-10, 
    8.868973e-10, 8.846992e-10, 8.835941e-10, 8.812664e-10, 8.816883e-10, 
    8.833963e-10, 8.872617e-10, 8.859469e-10, 8.892517e-10, 8.89177e-10, 
    8.928849e-10, 8.911984e-10, 8.97559e-10, 8.957414e-10, 9.009891e-10, 
    8.996703e-10, 9.009279e-10, 9.00546e-10, 9.009329e-10, 8.989984e-10, 
    8.998275e-10, 8.981237e-10, 8.915101e-10, 8.934425e-10, 8.877697e-10, 
    8.843905e-10, 8.82135e-10, 8.805373e-10, 8.807632e-10, 8.811946e-10, 
    8.834063e-10, 8.854818e-10, 8.870644e-10, 8.881235e-10, 8.891663e-10, 
    8.92343e-10, 8.940648e-10, 8.979287e-10, 8.972275e-10, 8.984124e-10, 
    8.995389e-10, 9.01435e-10, 9.011224e-10, 9.019586e-10, 8.983784e-10, 
    9.007593e-10, 8.968289e-10, 8.979046e-10, 8.894643e-10, 8.863009e-10, 
    8.849685e-10, 8.83791e-10, 8.809372e-10, 8.829089e-10, 8.82132e-10, 
    8.839772e-10, 8.851515e-10, 8.845701e-10, 8.881524e-10, 8.867604e-10, 
    8.94167e-10, 8.909383e-10, 8.994075e-10, 8.973711e-10, 8.99895e-10, 
    8.986065e-10, 9.008155e-10, 8.988273e-10, 9.022685e-10, 9.030193e-10, 
    9.025066e-10, 9.044711e-10, 8.987175e-10, 9.009294e-10, 8.845544e-10, 
    8.846494e-10, 8.850899e-10, 8.831538e-10, 8.830345e-10, 8.812556e-10, 
    8.828372e-10, 8.835118e-10, 8.852184e-10, 8.862304e-10, 8.871914e-10, 
    8.893037e-10, 8.916646e-10, 8.950578e-10, 8.975032e-10, 8.991433e-10, 
    8.981367e-10, 8.990255e-10, 8.980325e-10, 8.975664e-10, 9.027391e-10, 
    8.998362e-10, 9.041886e-10, 9.039473e-10, 9.01979e-10, 9.039745e-10, 
    8.847158e-10, 8.841701e-10, 8.822798e-10, 8.837591e-10, 8.810617e-10, 
    8.825735e-10, 8.834437e-10, 8.867927e-10, 8.875248e-10, 8.882082e-10, 
    8.895544e-10, 8.912835e-10, 8.943924e-10, 8.971177e-10, 8.996038e-10, 
    8.994214e-10, 8.994858e-10, 9.000427e-10, 8.986653e-10, 9.002686e-10, 
    9.005391e-10, 8.99834e-10, 9.039151e-10, 9.027492e-10, 9.039422e-10, 
    9.031827e-10, 8.843471e-10, 8.852646e-10, 8.847691e-10, 8.857017e-10, 
    8.850458e-10, 8.879661e-10, 8.888416e-10, 8.929623e-10, 8.912502e-10, 
    8.939862e-10, 8.915207e-10, 8.919473e-10, 8.940826e-10, 8.916496e-10, 
    8.969703e-10, 8.933597e-10, 9.000643e-10, 8.964636e-10, 9.002902e-10, 
    8.995931e-10, 9.007457e-10, 9.017795e-10, 9.030771e-10, 9.054751e-10, 
    9.049192e-10, 9.069218e-10, 8.86631e-10, 8.878221e-10, 8.877146e-10, 
    8.88959e-10, 8.898798e-10, 8.91872e-10, 8.9517e-10, 8.939269e-10, 
    8.962064e-10, 8.966653e-10, 8.932003e-10, 8.9533e-10, 8.886171e-10, 
    8.896877e-10, 8.890483e-10, 8.867265e-10, 8.942173e-10, 8.903413e-10, 
    8.975442e-10, 8.954124e-10, 9.016325e-10, 8.985424e-10, 9.046139e-10, 
    9.072152e-10, 9.096494e-10, 9.125082e-10, 8.884692e-10, 8.876602e-10, 
    8.891062e-10, 8.911114e-10, 8.929945e-10, 8.955429e-10, 8.958022e-10, 
    8.962808e-10, 8.975169e-10, 8.985576e-10, 8.964348e-10, 8.988182e-10, 
    8.899414e-10, 8.945573e-10, 8.873568e-10, 8.895049e-10, 8.90992e-10, 
    8.903369e-10, 8.937842e-10, 8.946108e-10, 8.979724e-10, 8.962326e-10, 
    9.065758e-10, 9.020018e-10, 9.146746e-10, 9.111374e-10, 8.873782e-10, 
    8.884651e-10, 8.922578e-10, 8.904493e-10, 8.957116e-10, 8.970219e-10, 
    8.980846e-10, 8.994474e-10, 8.995925e-10, 9.003994e-10, 8.990773e-10, 
    9.003462e-10, 8.955483e-10, 8.976921e-10, 8.918149e-10, 8.932413e-10, 
    8.925807e-10, 8.91864e-10, 8.940882e-10, 8.96469e-10, 8.965153e-10, 
    8.972799e-10, 8.994419e-10, 8.957329e-10, 9.071742e-10, 9.00118e-10, 
    8.896504e-10, 8.917493e-10, 8.920439e-10, 8.912317e-10, 8.968907e-10, 
    8.948307e-10, 9.003792e-10, 8.988787e-10, 9.013358e-10, 9.001153e-10, 
    8.99936e-10, 8.98367e-10, 8.973914e-10, 8.94926e-10, 8.929196e-10, 
    8.913489e-10, 8.917072e-10, 8.934465e-10, 8.966136e-10, 8.996076e-10, 
    8.989525e-10, 9.01149e-10, 8.953263e-10, 8.977705e-10, 8.968272e-10, 
    8.992857e-10, 8.938949e-10, 8.984991e-10, 8.9272e-10, 8.932257e-10, 
    8.947897e-10, 8.979393e-10, 8.986294e-10, 8.993745e-10, 8.989138e-10, 
    8.966932e-10, 8.963273e-10, 8.947507e-10, 8.943177e-10, 8.931152e-10, 
    8.921218e-10, 8.930306e-10, 8.939859e-10, 8.966923e-10, 8.991345e-10, 
    9.017949e-10, 9.02444e-10, 9.055623e-10, 9.030302e-10, 9.072144e-10, 
    9.036665e-10, 9.098022e-10, 8.987592e-10, 9.035531e-10, 8.948594e-10, 
    8.957946e-10, 8.974921e-10, 9.013747e-10, 8.992741e-10, 9.017285e-10, 
    8.963127e-10, 8.935092e-10, 8.927783e-10, 8.914435e-10, 8.928092e-10, 
    8.926964e-10, 8.940223e-10, 8.93596e-10, 8.967821e-10, 8.950701e-10, 
    8.999326e-10, 9.017079e-10, 9.067135e-10, 9.097832e-10, 9.12899e-10, 
    9.142764e-10, 9.146953e-10, 9.148706e-10,
  4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13,
  4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13,
  3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13,
  3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13,
  3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_UNSAT =
  0.6521466, 0.6199358, 0.6261668, 0.6004223, 0.6146694, 0.597862, 0.6455858, 
    0.6186643, 0.6358187, 0.6492325, 0.5513394, 0.5992808, 0.5029349, 
    0.5324775, 0.4592346, 0.5074909, 0.4498232, 0.4605904, 0.4285206, 
    0.4376057, 0.3977154, 0.4243563, 0.3777609, 0.4040047, 0.3998411, 
    0.4252484, 0.5895417, 0.557241, 0.5914716, 0.5868285, 0.5889112, 
    0.6143732, 0.6273103, 0.6546262, 0.6496472, 0.629595, 0.5847442, 
    0.5998703, 0.5619709, 0.5628186, 0.5215216, 0.5400124, 0.4719885, 
    0.4908208, 0.4372249, 0.4504615, 0.4378424, 0.4416528, 0.4377928, 
    0.4572741, 0.448883, 0.4661869, 0.5365321, 0.515565, 0.5789023, 
    0.6180338, 0.6443988, 0.6632628, 0.6605886, 0.6554966, 0.6294782, 
    0.6052585, 0.5869727, 0.5748302, 0.5629405, 0.5274277, 0.5089593, 
    0.4682146, 0.475395, 0.4632586, 0.4517877, 0.4328016, 0.4359025, 
    0.4276246, 0.4635788, 0.4395431, 0.4795039, 0.4684323, 0.5597121, 
    0.5957794, 0.611294, 0.6249675, 0.6585338, 0.635308, 0.6444404, 
    0.6227686, 0.6090942, 0.6158478, 0.5744992, 0.5904783, 0.507872, 
    0.5429558, 0.4531194, 0.4739178, 0.4481922, 0.461246, 0.4389758, 
    0.458998, 0.4245627, 0.4172216, 0.4222318, 0.4031411, 0.4601187, 
    0.4378416, 0.6160369, 0.614934, 0.6098035, 0.6324378, 0.6338297, 
    0.6547623, 0.6361294, 0.6282332, 0.6083047, 0.5965958, 0.5855246, 
    0.5613967, 0.5348251, 0.4984176, 0.4725581, 0.4557879, 0.4660424, 
    0.4569841, 0.4671147, 0.4718944, 0.4199648, 0.4488045, 0.4058613, 
    0.408186, 0.4274283, 0.4079238, 0.6141599, 0.6205116, 0.6426877, 
    0.6253165, 0.6570515, 0.6392404, 0.6290513, 0.590141, 0.5816863, 
    0.5738754, 0.5585446, 0.5390607, 0.5054522, 0.4765479, 0.4511244, 
    0.4529678, 0.4523183, 0.446711, 0.4606532, 0.4444395, 0.4417418, 
    0.448809, 0.4084978, 0.4198393, 0.4082355, 0.4156016, 0.6184453, 
    0.6077775, 0.6135358, 0.6027191, 0.6103334, 0.5766779, 0.5666953, 
    0.5207306, 0.5394415, 0.509775, 0.5364022, 0.5316489, 0.5088134, 
    0.5349518, 0.4780998, 0.5164932, 0.4464937, 0.4833831, 0.4442224, 
    0.4512331, 0.4396521, 0.4293905, 0.4166372, 0.3935757, 0.3988602, 
    0.3799428, 0.591968, 0.5783072, 0.5795079, 0.5653053, 0.5548706, 
    0.5324712, 0.4972155, 0.5103721, 0.4859704, 0.4812134, 0.5181221, 
    0.4955431, 0.5692184, 0.5570849, 0.5643007, 0.590886, 0.5073268, 
    0.5496942, 0.4721413, 0.4946553, 0.4308469, 0.4619408, 0.4017834, 
    0.3772648, 0.3549194, 0.3297415, 0.570893, 0.5801302, 0.5636239, 
    0.5410286, 0.520344, 0.4932884, 0.4901856, 0.485207, 0.472405, 0.4617463, 
    0.4836352, 0.4590902, 0.554279, 0.5037069, 0.5836322, 0.559163, 0.542353, 
    0.5497086, 0.5118842, 0.5031075, 0.4677585, 0.4856964, 0.3832431, 
    0.4272346, 0.3112941, 0.3416972, 0.5833675, 0.5709256, 0.5282783, 
    0.5484372, 0.4911327, 0.4775254, 0.4665761, 0.4527278, 0.4512443, 
    0.4431335, 0.4564569, 0.4436572, 0.4932313, 0.4706118, 0.5331001, 
    0.5177014, 0.5247661, 0.5325531, 0.508651, 0.4832871, 0.4827625, 
    0.4748749, 0.4529254, 0.4909075, 0.3777312, 0.4460846, 0.5574508, 
    0.5338964, 0.5305629, 0.5396284, 0.4788828, 0.5007936, 0.4433308, 
    0.458475, 0.4337767, 0.4459762, 0.4477833, 0.4636907, 0.4737087, 
    0.4997953, 0.5211511, 0.5383108, 0.5343038, 0.5155146, 0.4817786, 
    0.4511088, 0.4577561, 0.435633, 0.4955544, 0.4698261, 0.4795586, 
    0.4543518, 0.5107228, 0.462482, 0.5232685, 0.5178522, 0.5012258, 
    0.4681244, 0.4610138, 0.4534662, 0.4581179, 0.4809455, 0.4847285, 
    0.5016283, 0.5062345, 0.51903, 0.5297073, 0.5199482, 0.5097678, 
    0.4809369, 0.4558998, 0.4292449, 0.4228307, 0.3928166, 0.4171672, 
    0.3773654, 0.4110765, 0.3536533, 0.4597735, 0.4120944, 0.5004749, 
    0.4902615, 0.4727091, 0.4334483, 0.454469, 0.4299298, 0.4848772, 
    0.5148691, 0.522647, 0.5372615, 0.5223145, 0.5235248, 0.5093496, 0.51389, 
    0.4800051, 0.4982517, 0.447828, 0.4301219, 0.3819029, 0.3537589, 
    0.3263213, 0.3146154, 0.3111039, 0.3096431,
  0.9803318, 0.9605454, 0.9643664, 0.9485998, 0.9573179, 0.9470347, 
    0.9762947, 0.9597664, 0.9702914, 0.9785379, 0.9187019, 0.9479018, 
    0.8894453, 0.9072708, 0.8283049, 0.8921885, 0.8239651, 0.8289306, 
    0.8141972, 0.8183532, 0.8002158, 0.8122971, 0.7912525, 0.8030559, 
    0.8011748, 0.812704, 0.9419523, 0.9222851, 0.9431305, 0.9402968, 
    0.9415674, 0.9571369, 0.965069, 0.9818577, 0.978793, 0.9664704, 
    0.9390253, 0.9482616, 0.9251564, 0.9256718, 0.9006488, 0.9118317, 
    0.8342084, 0.8429748, 0.8181787, 0.8242584, 0.8184618, 0.8202091, 
    0.8184391, 0.827399, 0.8235319, 0.8315192, 0.9097244, 0.897054, 0.935463, 
    0.959381, 0.9755649, 0.9871783, 0.9855303, 0.9823941, 0.9663987, 
    0.9515567, 0.9403841, 0.9329814, 0.9257459, 0.904219, 0.8930725, 
    0.832459, 0.8357897, 0.8301644, 0.8248691, 0.816154, 0.8175731, 
    0.8137885, 0.8303121, 0.8192418, 0.8376997, 0.8325593, 0.9237867, 
    0.9457614, 0.9552522, 0.9636308, 0.9842645, 0.9699781, 0.9755906, 
    0.9622816, 0.953904, 0.9580396, 0.9327798, 0.9425239, 0.8924176, 
    0.9136155, 0.8254827, 0.8351038, 0.8232139, 0.8292333, 0.8189815, 
    0.8281947, 0.8123914, 0.8090492, 0.8113292, 0.8026649, 0.8287124, 
    0.8184617, 0.9581556, 0.95748, 0.954338, 0.9682155, 0.96907, 0.9819417, 
    0.9704822, 0.9656344, 0.9534206, 0.9462603, 0.9395008, 0.9248077, 
    0.9086917, 0.8867278, 0.8344727, 0.826713, 0.8314521, 0.8272649, 
    0.8319488, 0.8341644, 0.8102971, 0.823496, 0.8038954, 0.804948, 
    0.8136989, 0.8048292, 0.9570058, 0.9608977, 0.9745127, 0.9638444, 
    0.9833513, 0.9723939, 0.9661369, 0.9423187, 0.9371597, 0.9324002, 
    0.9230742, 0.9112552, 0.8909598, 0.8363258, 0.8245634, 0.8254126, 
    0.8251135, 0.8225328, 0.8289595, 0.8214888, 0.8202503, 0.8234978, 
    0.8050893, 0.8102396, 0.8049704, 0.8083124, 0.9596312, 0.9530981, 
    0.9566234, 0.9500037, 0.9546629, 0.934108, 0.9280307, 0.9001719, 
    0.9114861, 0.8935635, 0.9096456, 0.9067696, 0.8929855, 0.9087675, 
    0.8370477, 0.8976149, 0.8224329, 0.8395072, 0.8213891, 0.8246135, 
    0.8192913, 0.8145948, 0.8087832, 0.7983494, 0.8007315, 0.7922284, 
    0.9434334, 0.9351004, 0.9358316, 0.927184, 0.9208429, 0.9072666, 
    0.8860048, 0.8939226, 0.8407114, 0.8384954, 0.8985962, 0.8850001, 
    0.9295652, 0.9221885, 0.9265733, 0.9427732, 0.8920889, 0.9177018, 
    0.8342793, 0.8844663, 0.8152603, 0.8295553, 0.8020515, 0.7910313, 
    0.7810913, 0.7700264, 0.9305842, 0.9362109, 0.9261614, 0.9124481, 
    0.8999377, 0.8836454, 0.8426782, 0.8403557, 0.8344014, 0.8294646, 
    0.8396237, 0.8282372, 0.9204859, 0.8899093, 0.9383467, 0.9234512, 
    0.9132502, 0.9177098, 0.8948338, 0.8895479, 0.8322476, 0.8405837, 
    0.7937079, 0.813611, 0.7620181, 0.7752622, 0.9381848, 0.9306037, 
    0.9047318, 0.9169385, 0.8431205, 0.8367799, 0.8316993, 0.8253025, 
    0.8246188, 0.8208891, 0.8270217, 0.8211294, 0.8836111, 0.8335697, 
    0.907647, 0.8983426, 0.9026082, 0.907316, 0.8928856, 0.8394617, 
    0.8392166, 0.8355485, 0.825396, 0.8430154, 0.7912413, 0.8222472, 
    0.9224097, 0.90813, 0.9061126, 0.9115989, 0.8374111, 0.8881562, 
    0.8209796, 0.8279532, 0.8165999, 0.8221949, 0.8230259, 0.8303638, 
    0.8350067, 0.8875559, 0.9004251, 0.9108008, 0.9083753, 0.8970234, 
    0.8387591, 0.8245567, 0.8276218, 0.8174496, 0.8850064, 0.8332057, 
    0.8377258, 0.8260508, 0.8941342, 0.8298072, 0.9017034, 0.8984334, 
    0.8884161, 0.8324175, 0.829126, 0.8256428, 0.8277883, 0.8383711, 
    0.8401328, 0.888658, 0.8914307, 0.8991441, 0.9055949, 0.8996986, 
    0.893559, 0.8383668, 0.826765, 0.8145283, 0.8116018, 0.7980089, 
    0.8090253, 0.7910779, 0.8062613, 0.7805332, 0.8285543, 0.8067215, 
    0.8879642, 0.8427136, 0.8345433, 0.8164507, 0.8261049, 0.8148417, 
    0.840202, 0.8966346, 0.901328, 0.9101657, 0.9011273, 0.9018583, 
    0.8933064, 0.8960431, 0.8379331, 0.8866274, 0.8230467, 0.8149294, 
    0.7931064, 0.7805788, 0.7685341, 0.7634528, 0.7619358, 0.7613057,
  1.164523, 1.165765, 1.165546, 1.166379, 1.165941, 1.166451, 1.164798, 
    1.165808, 1.165187, 1.164647, 1.167402, 1.166411, 1.167567, 1.167575, 
    1.207638, 1.167592, 1.205625, 1.207926, 1.200946, 1.202963, 1.19385, 
    1.200011, 1.189015, 1.195333, 1.194353, 1.200212, 1.166672, 1.167321, 
    1.166623, 1.16674, 1.166688, 1.165951, 1.165505, 1.164417, 1.16463, 
    1.165421, 1.16679, 1.166395, 1.167248, 1.167235, 1.167614, 1.167522, 
    1.210318, 1.214179, 1.202879, 1.205762, 1.203015, 1.203851, 1.203004, 
    1.207221, 1.205422, 1.209106, 1.167549, 1.167614, 1.166924, 1.165829, 
    1.164847, 1.164034, 1.164154, 1.164379, 1.165426, 1.166237, 1.166736, 
    1.167011, 1.167233, 1.167598, 1.167598, 1.20953, 1.211025, 1.20849, 
    1.206048, 1.201901, 1.202587, 1.200746, 1.208557, 1.203389, 1.211872, 
    1.209576, 1.167284, 1.166508, 1.16605, 1.165589, 1.164246, 1.165206, 
    1.164845, 1.165667, 1.16612, 1.165903, 1.167017, 1.166648, 1.167594, 
    1.167495, 1.206334, 1.210719, 1.205273, 1.208064, 1.203264, 1.207588, 
    1.200058, 1.198392, 1.199531, 1.195131, 1.207826, 1.203015, 1.165896, 
    1.165933, 1.166097, 1.165316, 1.165263, 1.164411, 1.165175, 1.165471, 
    1.166144, 1.166486, 1.166771, 1.167258, 1.167561, 1.167534, 1.210436, 
    1.206904, 1.209075, 1.20716, 1.2093, 1.210298, 1.199017, 1.205405, 
    1.195768, 1.196309, 1.200702, 1.196248, 1.165958, 1.165745, 1.164916, 
    1.165577, 1.164311, 1.165053, 1.165441, 1.166657, 1.166862, 1.16703, 
    1.167302, 1.16753, 1.167582, 1.211263, 1.205905, 1.206301, 1.206162, 
    1.204952, 1.207939, 1.204459, 1.20387, 1.205406, 1.196382, 1.198988, 
    1.196321, 1.198021, 1.165816, 1.16616, 1.165978, 1.166312, 1.166081, 
    1.166972, 1.167167, 1.167614, 1.167527, 1.167601, 1.16755, 1.16758, 
    1.167597, 1.16756, 1.211583, 1.167615, 1.204905, 1.212667, 1.204412, 
    1.205928, 1.203413, 1.201141, 1.198258, 1.192863, 1.194121, 1.189554, 
    1.16661, 1.166937, 1.166911, 1.167192, 1.167356, 1.167575, 1.167524, 
    1.167603, 1.213195, 1.212223, 1.167616, 1.167508, 1.167121, 1.167324, 
    1.167209, 1.166638, 1.167591, 1.167422, 1.21035, 1.1675, 1.201466, 
    1.208211, 1.194812, 1.188892, 1.183216, 1.176446, 1.167089, 1.166897, 
    1.167221, 1.167513, 1.167615, 1.167485, 1.21405, 1.213039, 1.210404, 
    1.20817, 1.212719, 1.207608, 1.167363, 1.167572, 1.166816, 1.167293, 
    1.167501, 1.167422, 1.167608, 1.167569, 1.209435, 1.213139, 1.190364, 
    1.200658, 1.171193, 1.179714, 1.166823, 1.167089, 1.167595, 1.167437, 
    1.214242, 1.211465, 1.209187, 1.20625, 1.205931, 1.204174, 1.207047, 
    1.204288, 1.167485, 1.210031, 1.167572, 1.167616, 1.167607, 1.167575, 
    1.167597, 1.212647, 1.21254, 1.210917, 1.206292, 1.214196, 1.189008, 
    1.204816, 1.167319, 1.167567, 1.167585, 1.167525, 1.211744, 1.167553, 
    1.204217, 1.207477, 1.202117, 1.204793, 1.205184, 1.208581, 1.210675, 
    1.167545, 1.167614, 1.167536, 1.167564, 1.167614, 1.212339, 1.205902, 
    1.207324, 1.202528, 1.167508, 1.209867, 1.211883, 1.206598, 1.167604, 
    1.208326, 1.167611, 1.167616, 1.167556, 1.209512, 1.208015, 1.206408, 
    1.207401, 1.212168, 1.212942, 1.167559, 1.167586, 1.167616, 1.16759, 
    1.167615, 1.167601, 1.212166, 1.206928, 1.201108, 1.199667, 1.192682, 
    1.198379, 1.188917, 1.196979, 1.182886, 1.207752, 1.197214, 1.167551, 
    1.214066, 1.210467, 1.202044, 1.206623, 1.201261, 1.212972, 1.167613, 
    1.167612, 1.167544, 1.167613, 1.16761, 1.1676, 1.167612, 1.211975, 
    1.167533, 1.205194, 1.201304, 1.190036, 1.182914, 1.175492, 1.172158, 
    1.171137, 1.170709,
  0.5108873, 0.5006453, 0.5026345, 0.494389, 0.498961, 0.493565, 0.5088091, 
    0.5002388, 0.505708, 0.5099648, 0.4784437, 0.4940217, 0.4623524, 
    0.472223, 0.447545, 0.4638854, 0.4442539, 0.4480174, 0.4367121, 0.439945, 
    0.4255486, 0.4352217, 0.4181289, 0.427855, 0.4263298, 0.4355415, 
    0.4908817, 0.4803786, 0.4915048, 0.4900048, 0.490678, 0.4988661, 
    0.5029989, 0.5116718, 0.5100961, 0.5037271, 0.4893305, 0.4942116, 
    0.4819261, 0.482203, 0.4685815, 0.4747151, 0.4519686, 0.458429, 
    0.4398099, 0.444478, 0.4400288, 0.4413771, 0.4400112, 0.4468615, 
    0.4439239, 0.4499615, 0.4735652, 0.4665924, 0.4874378, 0.5000371, 
    0.5084326, 0.5144002, 0.5135561, 0.511947, 0.5036899, 0.4959436, 
    0.4900515, 0.4861158, 0.4822428, 0.4705471, 0.4643787, 0.4506639, 
    0.4531433, 0.4489452, 0.444943, 0.4382385, 0.4393408, 0.4363919, 
    0.4490565, 0.4406311, 0.4545566, 0.4507394, 0.4811872, 0.4928942, 
    0.4978797, 0.5022519, 0.512907, 0.5055455, 0.5084458, 0.5015501, 
    0.4971747, 0.4993382, 0.4860083, 0.4911842, 0.4640135, 0.475686, 
    0.4454094, 0.4526343, 0.4436812, 0.4482456, 0.4404303, 0.4474628, 
    0.4352957, 0.4326551, 0.4344591, 0.4275392, 0.4478532, 0.4400285, 
    0.4993987, 0.4990457, 0.4974021, 0.5046323, 0.5050753, 0.5117149, 
    0.5058067, 0.5032932, 0.4969214, 0.4931573, 0.4895831, 0.4817384, 
    0.4730004, 0.4608283, 0.4521652, 0.4463426, 0.4499115, 0.4467604, 
    0.4502831, 0.4519362, 0.4336439, 0.4438963, 0.428533, 0.4293803, 
    0.4363216, 0.4292848, 0.4987979, 0.5008293, 0.5078898, 0.5023633, 
    0.5124387, 0.5067953, 0.5035539, 0.4910752, 0.4883404, 0.4858055, 
    0.4808057, 0.4744009, 0.4632, 0.4535402, 0.4447105, 0.4453564, 0.4451289, 
    0.4431604, 0.4480393, 0.4423605, 0.4414085, 0.4438979, 0.4294938, 
    0.4335988, 0.4293983, 0.4320701, 0.500169, 0.4967523, 0.4985981, 
    0.4951277, 0.497572, 0.4867158, 0.4834679, 0.4683176, 0.4745266, 
    0.4646525, 0.4735223, 0.4719483, 0.4643295, 0.4730425, 0.4540739, 
    0.4669026, 0.4430839, 0.455887, 0.4422839, 0.4447486, 0.4406697, 
    0.4370227, 0.4324442, 0.4240225, 0.4259696, 0.4189483, 0.4916651, 
    0.4872447, 0.4876343, 0.4830147, 0.4796025, 0.4722209, 0.460422, 
    0.464853, 0.4567728, 0.4551434, 0.4674472, 0.4598562, 0.4842902, 
    0.4803277, 0.4826868, 0.4913158, 0.4638303, 0.4779036, 0.4520214, 
    0.4595557, 0.4375422, 0.4484872, 0.4270422, 0.4179423, 0.4094223, 
    0.3995158, 0.4848354, 0.4878361, 0.482466, 0.4750504, 0.4681888, 
    0.4590926, 0.4582124, 0.4565116, 0.4521125, 0.4484196, 0.4559734, 
    0.4474949, 0.4794082, 0.4626125, 0.4889706, 0.4810079, 0.4754873, 
    0.4779084, 0.46536, 0.4624107, 0.450506, 0.4566791, 0.4201835, 0.4362522, 
    0.3920159, 0.4042638, 0.488885, 0.4848461, 0.4708299, 0.4774906, 
    0.4585353, 0.4538765, 0.4500965, 0.4452723, 0.4447525, 0.4418998, 
    0.4465763, 0.4420846, 0.4590732, 0.4514931, 0.4724293, 0.4673066, 
    0.4696623, 0.4722481, 0.4642753, 0.4558541, 0.4556746, 0.4529641, 
    0.445341, 0.4584586, 0.4181173, 0.4429395, 0.4804477, 0.4726929, 
    0.4715882, 0.4745884, 0.4543432, 0.4616306, 0.4419695, 0.4472805, 
    0.4385855, 0.4429018, 0.4435375, 0.4490954, 0.4525622, 0.4612936, 
    0.468458, 0.4741532, 0.472828, 0.4665756, 0.4553371, 0.444705, 0.4470297, 
    0.4392451, 0.4598601, 0.4512215, 0.4545753, 0.4458406, 0.4649706, 
    0.448675, 0.4691637, 0.4673571, 0.4617764, 0.4506326, 0.4481648, 
    0.4455308, 0.447156, 0.4550514, 0.4563479, 0.4619121, 0.4634632, 
    0.4677504, 0.4713044, 0.4680568, 0.4646502, 0.4550485, 0.4463817, 
    0.4369707, 0.4346743, 0.4237417, 0.4326353, 0.4179798, 0.4304304, 
    0.4089319, 0.4477327, 0.4308, 0.4615231, 0.4582383, 0.4522173, 0.4384685, 
    0.4458816, 0.437215, 0.4563988, 0.4663596, 0.4689566, 0.4738064, 
    0.4688458, 0.469249, 0.4645099, 0.466032, 0.4547287, 0.4607723, 
    0.4435532, 0.4372836, 0.4196825, 0.4089731, 0.398142, 0.3933829, 
    0.3919375, 0.3913335,
  0.05040629, 0.04850325, 0.04886982, 0.04735983, 0.04819401, 0.0472103, 
    0.05001701, 0.04842853, 0.04943909, 0.05023329, 0.04451054, 0.04729316, 
    0.04172918, 0.04342415, 0.03924535, 0.04199011, 0.03870589, 0.03932309, 
    0.03748433, 0.03800546, 0.03571343, 0.03724534, 0.03456097, 0.03607566, 
    0.03583591, 0.03729654, 0.04672512, 0.04485133, 0.04683756, 0.04656712, 
    0.04668839, 0.04817662, 0.04893714, 0.05055368, 0.0502579, 0.0490718, 
    0.04644584, 0.04732761, 0.04512488, 0.04517392, 0.04279473, 0.0438577, 
    0.03997656, 0.04105711, 0.03798363, 0.0387425, 0.03801903, 0.03823752, 
    0.03801619, 0.039133, 0.03865201, 0.03964392, 0.04365737, 0.04245295, 
    0.04610626, 0.04839147, 0.04994667, 0.05106797, 0.05090855, 0.05060542, 
    0.04906491, 0.04764261, 0.04657554, 0.04586987, 0.04518098, 0.04313387, 
    0.04207425, 0.03976016, 0.04017192, 0.03947603, 0.03881852, 0.03772992, 
    0.03790778, 0.03743291, 0.03949441, 0.03811654, 0.04040762, 0.03977266, 
    0.04499416, 0.04708877, 0.04799602, 0.04879921, 0.05078616, 0.04940891, 
    0.04994912, 0.04866983, 0.04786717, 0.04826317, 0.04585067, 0.04677968, 
    0.04201196, 0.04402721, 0.03889485, 0.04008721, 0.03861242, 0.03936068, 
    0.03808402, 0.03923182, 0.03725718, 0.03683562, 0.03712336, 0.03602596, 
    0.03929606, 0.03801898, 0.04827427, 0.04820954, 0.04790872, 0.04923946, 
    0.04932162, 0.05056177, 0.04945744, 0.04899154, 0.04782094, 0.04713641, 
    0.04649125, 0.04509166, 0.04355915, 0.04147061, 0.04000923, 0.03904781, 
    0.03963565, 0.03911638, 0.03969712, 0.03997118, 0.03699318, 0.03864751, 
    0.03618252, 0.03631626, 0.03742164, 0.03630118, 0.04816412, 0.04853712, 
    0.04984533, 0.04881977, 0.05069794, 0.04964133, 0.04903974, 0.04676001, 
    0.04626804, 0.04581447, 0.04492676, 0.0438029, 0.04187335, 0.04023804, 
    0.0387805, 0.03888616, 0.03884894, 0.0385275, 0.0393267, 0.03839729, 
    0.03824261, 0.03864777, 0.03633419, 0.03698599, 0.03631911, 0.03674256, 
    0.0484157, 0.04779005, 0.04812751, 0.04749409, 0.04793976, 0.04597708, 
    0.04539829, 0.0427493, 0.04382483, 0.042121, 0.0436499, 0.04337651, 
    0.04206587, 0.04356647, 0.04032704, 0.04250616, 0.03851505, 0.04063014, 
    0.03838484, 0.03878673, 0.03812281, 0.03753423, 0.03680206, 0.0354748, 
    0.03577942, 0.03468728, 0.0468665, 0.04607169, 0.04614146, 0.04531783, 
    0.04471448, 0.0434238, 0.04140183, 0.04215525, 0.04077867, 0.04050568, 
    0.04259965, 0.04130614, 0.04554446, 0.04484237, 0.04525968, 0.04680343, 
    0.04198073, 0.04441566, 0.03998533, 0.04125536, 0.03761779, 0.03940049, 
    0.03594779, 0.03453223, 0.03323349, 0.03175559, 0.04564152, 0.04617761, 
    0.04522052, 0.04391619, 0.04272714, 0.04117716, 0.04102064, 0.04073485, 
    0.04000046, 0.03938936, 0.04064463, 0.0392371, 0.04468025, 0.0417734, 
    0.04638117, 0.04496247, 0.04399248, 0.04441652, 0.04224192, 0.0417391, 
    0.03973401, 0.04076294, 0.03487814, 0.0374105, 0.03065969, 0.0324596, 
    0.04636579, 0.04564342, 0.04318279, 0.04434318, 0.04107502, 0.04029411, 
    0.03966624, 0.0388724, 0.03878737, 0.03832241, 0.03908616, 0.03835244, 
    0.04117391, 0.03989763, 0.04345997, 0.0425755, 0.04298104, 0.04342851, 
    0.04205662, 0.04062465, 0.04059457, 0.04014208, 0.03888363, 0.0410621, 
    0.03455918, 0.03849152, 0.04486355, 0.04350572, 0.04331409, 0.0438356, 
    0.04037198, 0.04160662, 0.03833372, 0.03920184, 0.03778586, 0.03848539, 
    0.03858897, 0.03950083, 0.04007522, 0.04154947, 0.04277346, 0.04375975, 
    0.04352919, 0.04245006, 0.04053809, 0.0387796, 0.03916062, 0.03789233, 
    0.0413068, 0.03985256, 0.04041073, 0.03896549, 0.04217534, 0.03943145, 
    0.04289503, 0.04258417, 0.04163137, 0.03975498, 0.03934737, 0.03891472, 
    0.03918137, 0.0404903, 0.04070738, 0.04165441, 0.04191817, 0.04265175, 
    0.04326493, 0.04270443, 0.0421206, 0.04048982, 0.03905421, 0.03752587, 
    0.03715776, 0.03543098, 0.03683246, 0.03453799, 0.03648238, 0.03315951, 
    0.03927622, 0.03654094, 0.04158839, 0.04102501, 0.04001787, 0.03776699, 
    0.03897221, 0.03756515, 0.04071592, 0.04241303, 0.04285935, 0.04369935, 
    0.04284026, 0.04290975, 0.04209666, 0.04235691, 0.04043636, 0.04146114, 
    0.03859153, 0.03757618, 0.03480067, 0.03316571, 0.03155337, 0.03085798, 
    0.03064834, 0.03056096,
  0.001354541, 0.001276427, 0.00129135, 0.001230264, 0.001263885, 0.00122427, 
    0.001338433, 0.001273393, 0.001314641, 0.001347374, 0.001117798, 
    0.00122759, 0.001011639, 0.0010759, 0.0009199579, 0.001021442, 
    0.0009004449, 0.0009227818, 0.0008567956, 0.0008753256, 0.000794859, 
    0.0008483435, 0.0007559625, 0.000807397, 0.0007990908, 0.000850152, 
    0.001204892, 0.001131054, 0.001209373, 0.001198604, 0.001203429, 
    0.001263181, 0.001294097, 0.001360657, 0.001348393, 0.001299597, 
    0.001193785, 0.001228972, 0.001141734, 0.001143652, 0.001051878, 
    0.001092555, 0.000946636, 0.0009865368, 0.0008745463, 0.0009017646, 
    0.0008758098, 0.0008836208, 0.0008757084, 0.0009158821, 0.000898504, 
    0.0009344672, 0.001084848, 0.001038913, 0.001180328, 0.001271888, 
    0.001335529, 0.001382072, 0.001375421, 0.001362806, 0.001299316, 
    0.001241626, 0.001198939, 0.001170992, 0.001143928, 0.001064799, 
    0.001024611, 0.0009387132, 0.000953808, 0.000928346, 0.0009045069, 
    0.0008655111, 0.000871842, 0.0008549746, 0.0009290152, 0.000879293, 
    0.0009624854, 0.0009391702, 0.001136626, 0.001219406, 0.001255877, 
    0.00128847, 0.001370323, 0.001313403, 0.001335631, 0.001283201, 
    0.001250675, 0.001266686, 0.001170234, 0.001207066, 0.001022265, 
    0.00109909, 0.0009072636, 0.0009506955, 0.0008970787, 0.0009241484, 
    0.0008781307, 0.0009194668, 0.0008487616, 0.0008339213, 0.0008440409, 
    0.0008056728, 0.0009217996, 0.0008758079, 0.001267136, 0.001264513, 
    0.001252351, 0.001306457, 0.001309823, 0.001360993, 0.001315395, 
    0.001296318, 0.00124881, 0.001221312, 0.001195589, 0.001140435, 
    0.001081077, 0.001001956, 0.0009478338, 0.0009127961, 0.0009341651, 
    0.0009152799, 0.0009364096, 0.0009464385, 0.0008394574, 0.0008983418, 
    0.0008111087, 0.0008157624, 0.0008545757, 0.0008152371, 0.001262675, 
    0.001277803, 0.00133135, 0.001289308, 0.001366652, 0.00132295, 
    0.001298287, 0.001206282, 0.001186733, 0.001168807, 0.001133996, 
    0.001090445, 0.001017052, 0.0009562392, 0.0009031352, 0.0009069498, 
    0.0009056053, 0.0008940244, 0.000922913, 0.0008893474, 0.000883803, 
    0.0008983515, 0.0008163871, 0.0008392044, 0.0008158616, 0.0008306575, 
    0.001272872, 0.001247565, 0.001261193, 0.001235654, 0.001253605, 
    0.001175223, 0.001152442, 0.001050152, 0.001091289, 0.001026373, 
    0.001084562, 0.001074076, 0.001024295, 0.001081358, 0.0009595156, 
    0.001040927, 0.0008935765, 0.0009707024, 0.0008889008, 0.00090336, 
    0.0008795169, 0.0008585642, 0.0008327438, 0.0007866363, 0.000797138, 
    0.0007597107, 0.001210527, 0.001178961, 0.001181721, 0.001149287, 
    0.001125725, 0.001075887, 0.0009993853, 0.001027664, 0.0009762007, 
    0.0009661037, 0.001044471, 0.0009958127, 0.001158181, 0.001130705, 
    0.001147009, 0.001208012, 0.001021089, 0.001114118, 0.0009469572, 
    0.000993919, 0.0008615279, 0.0009255962, 0.0008029632, 0.0007549848, 
    0.0007112785, 0.00066267, 0.001161997, 0.001183152, 0.001145476, 
    0.001094808, 0.00104931, 0.0009910051, 0.000985181, 0.0009745774, 
    0.0009475121, 0.0009251914, 0.0009712384, 0.0009196587, 0.001124393, 
    0.001013298, 0.001191218, 0.001135389, 0.00109775, 0.001114151, 
    0.001030935, 0.001012011, 0.0009377576, 0.0009756181, 0.0007662062, 
    0.0008541814, 0.0006274168, 0.0006856739, 0.001190608, 0.001162071, 
    0.001066667, 0.001111309, 0.000987203, 0.000958303, 0.000935282, 
    0.0009064524, 0.0009033831, 0.0008866618, 0.0009141851, 0.0008877386, 
    0.0009908836, 0.0009437434, 0.001077273, 0.001043555, 0.00105897, 
    0.001076067, 0.001023947, 0.0009704994, 0.0009693875, 0.0009527111, 
    0.0009068582, 0.0009867223, 0.0007559014, 0.000892731, 0.001131531, 
    0.001079027, 0.001071687, 0.001091704, 0.0009611713, 0.001007045, 
    0.0008870675, 0.0009183789, 0.0008675006, 0.0008925106, 0.0008962351, 
    0.000929249, 0.0009502553, 0.001004905, 0.00105107, 0.001088784, 
    0.001079928, 0.001038803, 0.0009673006, 0.0009031026, 0.0009168835, 
    0.0008712913, 0.0009958376, 0.0009420934, 0.0009626002, 0.0009098172, 
    0.001028422, 0.0009267227, 0.001055694, 0.001043884, 0.001007972, 
    0.0009385237, 0.0009236644, 0.0009079817, 0.0009176364, 0.0009655358, 
    0.0009735606, 0.001008835, 0.001018736, 0.001046447, 0.001069806, 
    0.001048447, 0.001026358, 0.000965518, 0.0009130279, 0.0008582677, 
    0.0008452535, 0.0007851294, 0.0008338104, 0.0007551809, 0.0008215553, 
    0.0007088166, 0.000921079, 0.000823601, 0.001006362, 0.000985343, 
    0.0009481506, 0.0008668292, 0.0009100602, 0.0008596604, 0.0009738766, 
    0.001037402, 0.001054336, 0.001086462, 0.00105361, 0.001056254, 
    0.001025455, 0.001035279, 0.0009635453, 0.001001601, 0.0008963271, 
    0.0008600517, 0.0007635673, 0.000709023, 0.000656114, 0.0006337448, 
    0.0006270551, 0.0006242744,
  8.907522e-06, 8.124075e-06, 8.271948e-06, 7.672142e-06, 8.000457e-06, 
    7.614084e-06, 8.744086e-06, 8.094111e-06, 8.504462e-06, 8.834687e-06, 
    6.607358e-06, 7.646223e-06, 5.652549e-06, 6.224463e-06, 4.870591e-06, 
    5.738567e-06, 4.709587e-06, 4.894054e-06, 4.356659e-06, 4.505246e-06, 
    3.873723e-06, 4.2895e-06, 3.2485e-06, 3.969741e-06, 3.906031e-06, 
    4.303837e-06, 7.427361e-06, 6.730098e-06, 7.470406e-06, 7.367106e-06, 
    7.413332e-06, 7.993537e-06, 8.299263e-06, 8.969827e-06, 8.845029e-06, 
    8.354045e-06, 7.321032e-06, 7.65961e-06, 6.829527e-06, 6.847439e-06, 
    6.008459e-06, 6.375738e-06, 5.093856e-06, 5.43438e-06, 4.498961e-06, 
    4.720414e-06, 4.509154e-06, 4.572358e-06, 4.508336e-06, 4.8368e-06, 
    4.69368e-06, 4.991572e-06, 6.305586e-06, 5.892961e-06, 7.192882e-06, 
    8.07927e-06, 8.714725e-06, 9.189076e-06, 9.120808e-06, 8.991758e-06, 
    8.351236e-06, 7.782598e-06, 7.370309e-06, 7.104409e-06, 6.850017e-06, 
    6.124314e-06, 5.766464e-06, 5.027177e-06, 5.154486e-06, 4.940403e-06, 
    4.742942e-06, 4.426317e-06, 4.477172e-06, 4.342156e-06, 4.945987e-06, 
    4.537299e-06, 5.228183e-06, 5.031015e-06, 6.781909e-06, 7.567072e-06, 
    7.921852e-06, 8.243349e-06, 9.068585e-06, 8.492048e-06, 8.71575e-06, 
    8.191092e-06, 7.870924e-06, 8.028016e-06, 7.097248e-06, 7.448234e-06, 
    5.745803e-06, 6.435436e-06, 4.765626e-06, 5.128144e-06, 4.682011e-06, 
    4.905422e-06, 4.5279e-06, 4.866515e-06, 4.292813e-06, 4.175808e-06, 
    4.255462e-06, 3.956484e-06, 4.885888e-06, 4.509139e-06, 8.032442e-06, 
    8.006639e-06, 7.887328e-06, 8.422528e-06, 8.456195e-06, 8.973255e-06, 
    8.512015e-06, 8.32137e-06, 7.852695e-06, 7.585482e-06, 7.338266e-06, 
    6.817408e-06, 6.271351e-06, 5.568034e-06, 5.103964e-06, 4.811271e-06, 
    4.989043e-06, 4.831814e-06, 5.007849e-06, 5.09219e-06, 4.219315e-06, 
    4.692352e-06, 3.998338e-06, 4.034304e-06, 4.338982e-06, 4.030238e-06, 
    7.988565e-06, 8.137677e-06, 8.672525e-06, 8.251671e-06, 9.03104e-06, 
    8.587904e-06, 8.340985e-06, 7.440705e-06, 7.25378e-06, 7.083759e-06, 
    6.757432e-06, 6.356506e-06, 5.699986e-06, 5.175098e-06, 4.731668e-06, 
    4.763041e-06, 4.751975e-06, 4.657042e-06, 4.895144e-06, 4.618902e-06, 
    4.573837e-06, 4.692431e-06, 4.039141e-06, 4.217322e-06, 4.035072e-06, 
    4.150239e-06, 8.088973e-06, 7.840531e-06, 7.974009e-06, 7.724476e-06, 
    7.899594e-06, 7.144458e-06, 6.929709e-06, 5.993034e-06, 6.364196e-06, 
    5.781997e-06, 6.30298e-06, 6.207965e-06, 5.76368e-06, 6.273896e-06, 
    5.202919e-06, 5.91086e-06, 4.653385e-06, 5.298312e-06, 4.615265e-06, 
    4.733515e-06, 4.539111e-06, 4.370761e-06, 4.166577e-06, 3.811246e-06, 
    3.89111e-06, 3.609434e-06, 7.481508e-06, 7.179908e-06, 7.206108e-06, 
    6.900146e-06, 6.68066e-06, 6.224341e-06, 5.545674e-06, 5.793388e-06, 
    5.345422e-06, 5.259024e-06, 5.942381e-06, 5.51465e-06, 6.983602e-06, 
    6.726852e-06, 6.878819e-06, 7.457327e-06, 5.735462e-06, 6.573413e-06, 
    5.096567e-06, 5.498228e-06, 4.394431e-06, 4.917477e-06, 3.935684e-06, 
    3.243093e-06, 3.002658e-06, 2.738317e-06, 7.019516e-06, 7.219707e-06, 
    6.86448e-06, 6.396302e-06, 5.985518e-06, 5.472994e-06, 5.422681e-06, 
    5.331498e-06, 5.101249e-06, 4.914106e-06, 5.302898e-06, 4.868108e-06, 
    6.668323e-06, 5.667075e-06, 7.296533e-06, 6.770397e-06, 6.42318e-06, 
    6.573718e-06, 5.822279e-06, 5.655806e-06, 5.019156e-06, 5.340423e-06, 
    3.657726e-06, 4.335845e-06, 2.548767e-06, 2.862999e-06, 7.290711e-06, 
    7.02022e-06, 6.141126e-06, 6.547546e-06, 5.440129e-06, 5.192617e-06, 
    4.998398e-06, 4.758946e-06, 4.733705e-06, 4.597053e-06, 4.822754e-06, 
    4.605808e-06, 5.471943e-06, 5.069476e-06, 6.236884e-06, 5.93423e-06, 
    6.071952e-06, 6.225975e-06, 5.760613e-06, 5.296576e-06, 5.287068e-06, 
    5.145197e-06, 4.762287e-06, 5.43598e-06, 3.248162e-06, 4.646483e-06, 
    6.734522e-06, 6.252769e-06, 6.186384e-06, 6.367977e-06, 5.217e-06, 
    5.612399e-06, 4.600351e-06, 4.85749e-06, 4.442274e-06, 4.644685e-06, 
    4.67511e-06, 4.947939e-06, 5.124421e-06, 5.593733e-06, 6.001236e-06, 
    6.341383e-06, 6.260929e-06, 5.89199e-06, 5.269239e-06, 4.7314e-06, 
    4.845094e-06, 4.472739e-06, 5.514866e-06, 5.055587e-06, 5.229162e-06, 
    4.786674e-06, 5.800079e-06, 4.926864e-06, 6.042595e-06, 5.937155e-06, 
    5.620492e-06, 5.025586e-06, 4.901395e-06, 4.771541e-06, 4.851334e-06, 
    5.254179e-06, 5.322783e-06, 5.628036e-06, 5.714779e-06, 5.959987e-06, 
    6.169415e-06, 5.977821e-06, 5.781862e-06, 5.254027e-06, 4.813186e-06, 
    4.368395e-06, 4.265044e-06, 3.799838e-06, 4.174938e-06, 3.244177e-06, 
    4.079244e-06, 2.98919e-06, 4.879901e-06, 4.09516e-06, 5.60644e-06, 
    5.424079e-06, 5.106639e-06, 4.436887e-06, 4.788679e-06, 4.37951e-06, 
    5.325491e-06, 5.879554e-06, 6.030437e-06, 6.320253e-06, 6.023941e-06, 
    6.047612e-06, 5.773906e-06, 5.860736e-06, 5.237212e-06, 5.564952e-06, 
    4.675862e-06, 4.382634e-06, 3.638076e-06, 2.990319e-06, 2.702924e-06, 
    2.582651e-06, 2.546832e-06, 2.531964e-06,
  8.171993e-09, 6.97288e-09, 7.196179e-09, 6.299845e-09, 6.787349e-09, 
    6.214455e-09, 7.918667e-09, 6.927812e-09, 7.55021e-09, 8.0589e-09, 
    4.776885e-09, 6.261693e-09, 3.501304e-09, 4.253917e-09, 2.537115e-09, 
    3.612148e-09, 2.349385e-09, 2.564806e-09, 1.95272e-09, 2.117128e-09, 
    1.447282e-09, 1.879712e-09, 1.159808e-09, 1.544e-09, 1.479603e-09, 
    1.895228e-09, 5.941564e-09, 4.947489e-09, 6.004236e-09, 5.854079e-09, 
    5.921168e-09, 6.776995e-09, 7.237586e-09, 8.268986e-09, 8.074939e-09, 
    7.32078e-09, 5.787375e-09, 6.281392e-09, 5.086697e-09, 5.111869e-09, 
    3.965441e-09, 4.458813e-09, 2.8039e-09, 3.224183e-09, 2.110095e-09, 
    2.361882e-09, 2.121504e-09, 2.192643e-09, 2.120587e-09, 2.497382e-09, 
    2.331059e-09, 2.680776e-09, 4.363508e-09, 3.813253e-09, 5.602746e-09, 
    6.905513e-09, 7.87333e-09, 8.612099e-09, 8.504966e-09, 8.30318e-09, 
    7.31651e-09, 6.462988e-09, 5.858721e-09, 5.476063e-09, 5.115495e-09, 
    4.119555e-09, 3.648282e-09, 2.723465e-09, 2.877584e-09, 2.619748e-09, 
    2.387943e-09, 2.029309e-09, 2.085767e-09, 1.936884e-09, 2.626391e-09, 
    2.153098e-09, 2.967831e-09, 2.728078e-09, 5.019918e-09, 6.145498e-09, 
    6.669927e-09, 7.152878e-09, 8.423194e-09, 7.53122e-09, 7.874911e-09, 
    7.073898e-09, 6.594086e-09, 6.82862e-09, 5.465838e-09, 5.971936e-09, 
    3.621512e-09, 4.540297e-09, 2.414267e-09, 2.845506e-09, 2.317642e-09, 
    2.578253e-09, 2.142532e-09, 2.532314e-09, 1.883294e-09, 1.758042e-09, 
    1.843029e-09, 1.530528e-09, 2.555159e-09, 2.121487e-09, 6.835251e-09, 
    6.796603e-09, 6.618496e-09, 7.425056e-09, 7.47643e-09, 8.274328e-09, 
    7.56177e-09, 7.271135e-09, 6.566984e-09, 6.172482e-09, 5.812306e-09, 
    5.069683e-09, 4.317177e-09, 3.393258e-09, 2.816149e-09, 2.46748e-09, 
    2.67775e-09, 2.491534e-09, 2.700268e-09, 2.801883e-09, 1.80431e-09, 
    2.329531e-09, 1.573185e-09, 1.610132e-09, 1.933423e-09, 1.605942e-09, 
    6.769557e-09, 6.993357e-09, 7.808257e-09, 7.165472e-09, 8.3645e-09, 
    7.678108e-09, 7.300928e-09, 5.960976e-09, 5.690318e-09, 5.446589e-09, 
    4.985671e-09, 4.432636e-09, 3.562324e-09, 2.902749e-09, 2.374892e-09, 
    2.411264e-09, 2.398417e-09, 2.289004e-09, 2.566094e-09, 2.245458e-09, 
    2.194314e-09, 2.329622e-09, 1.615122e-09, 1.802184e-09, 1.610924e-09, 
    1.731022e-09, 6.92009e-09, 6.548912e-09, 6.747793e-09, 6.37703e-09, 
    6.63676e-09, 5.533328e-09, 5.227848e-09, 3.945032e-09, 4.443097e-09, 
    3.668441e-09, 4.359976e-09, 4.231711e-09, 3.644672e-09, 4.320618e-09, 
    2.936809e-09, 3.83674e-09, 2.284818e-09, 3.05439e-09, 2.241319e-09, 
    2.377028e-09, 2.155137e-09, 1.968154e-09, 1.748272e-09, 1.385431e-09, 
    1.464647e-09, 1.191778e-09, 6.020423e-09, 5.584127e-09, 5.62174e-09, 
    5.186104e-09, 4.878605e-09, 4.253753e-09, 3.364818e-09, 3.683243e-09, 
    3.112905e-09, 3.005816e-09, 3.878192e-09, 3.325459e-09, 5.304142e-09, 
    4.942961e-09, 5.156036e-09, 5.985178e-09, 3.608131e-09, 4.72995e-09, 
    2.807183e-09, 3.304675e-09, 1.994142e-09, 2.592532e-09, 1.509468e-09, 
    1.153147e-09, 8.742305e-10, 6.085717e-10, 5.355123e-09, 5.641283e-09, 
    5.135844e-09, 4.486841e-09, 3.935096e-09, 3.272802e-09, 3.209491e-09, 
    3.09558e-09, 2.812858e-09, 2.588537e-09, 3.060074e-09, 2.534189e-09, 
    4.861451e-09, 3.519961e-09, 5.751976e-09, 5.003804e-09, 4.52354e-09, 
    4.730371e-09, 3.720849e-09, 3.505485e-09, 2.713832e-09, 3.106682e-09, 
    1.237238e-09, 1.930005e-09, 4.463161e-10, 7.283275e-10, 5.743571e-09, 
    5.356122e-09, 4.142038e-09, 4.694256e-09, 3.231411e-09, 2.924184e-09, 
    2.688945e-09, 2.406508e-09, 2.377248e-09, 2.22062e-09, 2.480918e-09, 
    2.230564e-09, 3.271476e-09, 2.774416e-09, 4.270654e-09, 3.867463e-09, 
    4.049724e-09, 4.255953e-09, 3.640696e-09, 3.052239e-09, 3.040468e-09, 
    2.866261e-09, 2.410387e-09, 3.226194e-09, 1.159391e-09, 2.276924e-09, 
    4.953665e-09, 4.29208e-09, 4.202707e-09, 4.448244e-09, 2.954088e-09, 
    3.449869e-09, 2.224364e-09, 2.52169e-09, 2.046976e-09, 2.27487e-09, 
    2.309716e-09, 2.628713e-09, 2.840981e-09, 3.426021e-09, 3.955882e-09, 
    4.412078e-09, 4.303097e-09, 3.811979e-09, 3.018426e-09, 2.374581e-09, 
    2.507119e-09, 2.080828e-09, 3.325733e-09, 2.757658e-09, 2.969033e-09, 
    2.438765e-09, 3.691943e-09, 2.603666e-09, 4.010702e-09, 3.871313e-09, 
    3.460221e-09, 2.721553e-09, 2.573487e-09, 2.421144e-09, 2.51445e-09, 
    2.99984e-09, 3.084749e-09, 3.469877e-09, 3.581408e-09, 3.901393e-09, 
    4.179936e-09, 3.924928e-09, 3.668267e-09, 2.999653e-09, 2.46972e-09, 
    1.965563e-09, 1.853333e-09, 1.374232e-09, 1.75712e-09, 1.154481e-09, 
    1.656671e-09, 8.596314e-10, 2.548093e-09, 1.673252e-09, 3.442251e-09, 
    3.211246e-09, 2.819392e-09, 2.041006e-09, 2.441102e-09, 1.977749e-09, 
    3.088113e-09, 3.795681e-09, 3.994568e-09, 4.383393e-09, 3.985953e-09, 
    4.017364e-09, 3.657937e-09, 3.771054e-09, 2.978937e-09, 3.389335e-09, 
    2.31058e-09, 1.981178e-09, 1.218672e-09, 8.608512e-10, 5.764348e-10, 
    4.735223e-10, 4.447864e-10, 4.331205e-10,
  4.330855e-13, 4.283784e-13, 4.292556e-13, 4.257326e-13, 4.276493e-13, 
    4.253967e-13, 4.320918e-13, 4.282013e-13, 4.306457e-13, 4.326419e-13, 
    4.197344e-13, 4.255825e-13, 4.146965e-13, 4.176706e-13, 4.108788e-13, 
    4.151349e-13, 4.101342e-13, 4.109886e-13, 4.085595e-13, 4.092125e-13, 
    4.065496e-13, 4.082694e-13, 4.0541e-13, 4.069345e-13, 4.066782e-13, 
    4.083311e-13, 4.24323e-13, 4.204071e-13, 4.245696e-13, 4.239786e-13, 
    4.242427e-13, 4.276086e-13, 4.294182e-13, 4.33466e-13, 4.327048e-13, 
    4.297449e-13, 4.23716e-13, 4.2566e-13, 4.209559e-13, 4.210552e-13, 
    4.165313e-13, 4.184795e-13, 4.119361e-13, 4.136002e-13, 4.091845e-13, 
    4.101838e-13, 4.092298e-13, 4.095122e-13, 4.092262e-13, 4.107212e-13, 
    4.100615e-13, 4.114482e-13, 4.181033e-13, 4.159299e-13, 4.229891e-13, 
    4.281137e-13, 4.319139e-13, 4.348112e-13, 4.343912e-13, 4.336e-13, 
    4.297281e-13, 4.263742e-13, 4.239969e-13, 4.224902e-13, 4.210695e-13, 
    4.1714e-13, 4.152777e-13, 4.116174e-13, 4.12228e-13, 4.112064e-13, 
    4.102872e-13, 4.088637e-13, 4.090879e-13, 4.084966e-13, 4.112327e-13, 
    4.093552e-13, 4.125854e-13, 4.116357e-13, 4.206927e-13, 4.251254e-13, 
    4.271878e-13, 4.290855e-13, 4.340706e-13, 4.305712e-13, 4.319201e-13, 
    4.287752e-13, 4.268896e-13, 4.278115e-13, 4.224499e-13, 4.244425e-13, 
    4.151719e-13, 4.18801e-13, 4.103916e-13, 4.121009e-13, 4.100083e-13, 
    4.110419e-13, 4.093133e-13, 4.108597e-13, 4.082836e-13, 4.077858e-13, 
    4.081236e-13, 4.068809e-13, 4.109503e-13, 4.092298e-13, 4.278376e-13, 
    4.276857e-13, 4.269856e-13, 4.301544e-13, 4.303561e-13, 4.334869e-13, 
    4.306911e-13, 4.2955e-13, 4.267831e-13, 4.252316e-13, 4.238142e-13, 
    4.208889e-13, 4.179204e-13, 4.142691e-13, 4.119847e-13, 4.106026e-13, 
    4.114363e-13, 4.106981e-13, 4.115255e-13, 4.119281e-13, 4.079697e-13, 
    4.100555e-13, 4.070506e-13, 4.071976e-13, 4.084828e-13, 4.07181e-13, 
    4.275794e-13, 4.284588e-13, 4.316585e-13, 4.291349e-13, 4.338405e-13, 
    4.311478e-13, 4.296669e-13, 4.243993e-13, 4.233339e-13, 4.223741e-13, 
    4.205577e-13, 4.183762e-13, 4.149378e-13, 4.123277e-13, 4.102354e-13, 
    4.103797e-13, 4.103287e-13, 4.098947e-13, 4.109937e-13, 4.097218e-13, 
    4.095189e-13, 4.100558e-13, 4.072175e-13, 4.079613e-13, 4.072008e-13, 
    4.076784e-13, 4.281709e-13, 4.26712e-13, 4.274938e-13, 4.260362e-13, 
    4.270574e-13, 4.227157e-13, 4.215122e-13, 4.164506e-13, 4.184174e-13, 
    4.153574e-13, 4.180894e-13, 4.17583e-13, 4.152635e-13, 4.17934e-13, 
    4.124626e-13, 4.160227e-13, 4.098781e-13, 4.129281e-13, 4.097054e-13, 
    4.102439e-13, 4.093634e-13, 4.086208e-13, 4.07747e-13, 4.063034e-13, 
    4.066187e-13, 4.05532e-13, 4.246333e-13, 4.229158e-13, 4.230639e-13, 
    4.213477e-13, 4.201356e-13, 4.1767e-13, 4.141566e-13, 4.15416e-13, 
    4.131598e-13, 4.127358e-13, 4.161865e-13, 4.140009e-13, 4.218129e-13, 
    4.203893e-13, 4.212292e-13, 4.244946e-13, 4.15119e-13, 4.195493e-13, 
    4.119491e-13, 4.139186e-13, 4.087241e-13, 4.110985e-13, 4.067971e-13, 
    4.053835e-13, 4.042697e-13, 4.032074e-13, 4.220137e-13, 4.231409e-13, 
    4.211497e-13, 4.185901e-13, 4.164114e-13, 4.137925e-13, 4.13542e-13, 
    4.130912e-13, 4.119716e-13, 4.110827e-13, 4.129506e-13, 4.108672e-13, 
    4.200679e-13, 4.147703e-13, 4.235767e-13, 4.206292e-13, 4.187349e-13, 
    4.195509e-13, 4.155646e-13, 4.147131e-13, 4.115792e-13, 4.131351e-13, 
    4.057131e-13, 4.084693e-13, 4.025578e-13, 4.036865e-13, 4.235436e-13, 
    4.220177e-13, 4.172288e-13, 4.194085e-13, 4.136288e-13, 4.124126e-13, 
    4.114806e-13, 4.103608e-13, 4.102448e-13, 4.096233e-13, 4.106559e-13, 
    4.096628e-13, 4.137873e-13, 4.118193e-13, 4.177367e-13, 4.161441e-13, 
    4.168642e-13, 4.176787e-13, 4.152478e-13, 4.129196e-13, 4.12873e-13, 
    4.121831e-13, 4.103762e-13, 4.136081e-13, 4.054084e-13, 4.098467e-13, 
    4.204315e-13, 4.178213e-13, 4.174684e-13, 4.184377e-13, 4.12531e-13, 
    4.144931e-13, 4.096381e-13, 4.108176e-13, 4.089339e-13, 4.098386e-13, 
    4.099768e-13, 4.112419e-13, 4.12083e-13, 4.143987e-13, 4.164935e-13, 
    4.18295e-13, 4.178648e-13, 4.159248e-13, 4.127857e-13, 4.102342e-13, 
    4.107598e-13, 4.090683e-13, 4.140019e-13, 4.117529e-13, 4.125902e-13, 
    4.104888e-13, 4.154504e-13, 4.111426e-13, 4.167101e-13, 4.161593e-13, 
    4.14534e-13, 4.116098e-13, 4.11023e-13, 4.104189e-13, 4.107889e-13, 
    4.127122e-13, 4.130483e-13, 4.145722e-13, 4.150133e-13, 4.162782e-13, 
    4.173785e-13, 4.163712e-13, 4.153567e-13, 4.127114e-13, 4.106115e-13, 
    4.086105e-13, 4.081646e-13, 4.062588e-13, 4.077822e-13, 4.053888e-13, 
    4.073827e-13, 4.042114e-13, 4.109223e-13, 4.074487e-13, 4.144629e-13, 
    4.13549e-13, 4.119975e-13, 4.089102e-13, 4.104981e-13, 4.086589e-13, 
    4.130616e-13, 4.158604e-13, 4.166463e-13, 4.181818e-13, 4.166123e-13, 
    4.167364e-13, 4.153159e-13, 4.157631e-13, 4.126294e-13, 4.142536e-13, 
    4.099803e-13, 4.086726e-13, 4.056391e-13, 4.042163e-13, 4.030788e-13, 
    4.026668e-13, 4.025517e-13, 4.02505e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC =
  8.949655e-07, 8.949654e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949655e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 
    8.949653e-07, 8.949654e-07, 8.949652e-07, 8.949653e-07, 8.949651e-07, 
    8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.94965e-07, 8.949651e-07, 8.94965e-07, 8.949651e-07, 8.94965e-07, 
    8.949651e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949652e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 8.949654e-07, 
    8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949652e-07, 
    8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949652e-07, 8.949653e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.94965e-07, 8.949651e-07, 8.949651e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949652e-07, 8.949653e-07, 
    8.949652e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949653e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.94965e-07, 
    8.94965e-07, 8.94965e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949652e-07, 8.949653e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 8.94965e-07, 
    8.94965e-07, 8.94965e-07, 8.949649e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949652e-07, 8.949651e-07, 
    8.949653e-07, 8.949652e-07, 8.949654e-07, 8.949654e-07, 8.949653e-07, 
    8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.94965e-07, 8.949651e-07, 8.949648e-07, 8.949649e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949652e-07, 8.94965e-07, 8.949651e-07, 
    8.949654e-07, 8.949653e-07, 8.949653e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949653e-07, 8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949651e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949653e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949651e-07, 
    8.949651e-07, 8.949651e-07, 8.94965e-07, 8.949651e-07, 8.94965e-07, 
    8.949651e-07, 8.94965e-07, 8.949651e-07, 8.949651e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 8.949652e-07, 
    8.949651e-07, 8.949651e-07, 8.94965e-07, 8.94965e-07, 8.949649e-07, 
    8.949648e-07, 8.949648e-07, 8.949648e-07 ;

 CWDC_HR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC_LOSS =
  6.01737e-16, 6.033623e-16, 6.030466e-16, 6.043563e-16, 6.036301e-16, 
    6.044873e-16, 6.020669e-16, 6.034266e-16, 6.025589e-16, 6.018837e-16, 
    6.068941e-16, 6.044148e-16, 6.094675e-16, 6.07889e-16, 6.118515e-16, 
    6.092216e-16, 6.123814e-16, 6.117762e-16, 6.135982e-16, 6.130765e-16, 
    6.154034e-16, 6.13839e-16, 6.166091e-16, 6.150302e-16, 6.152771e-16, 
    6.137872e-16, 6.049145e-16, 6.065855e-16, 6.048154e-16, 6.050538e-16, 
    6.049469e-16, 6.03645e-16, 6.029881e-16, 6.016131e-16, 6.018629e-16, 
    6.028729e-16, 6.05161e-16, 6.04385e-16, 6.06341e-16, 6.062969e-16, 
    6.084711e-16, 6.074912e-16, 6.111412e-16, 6.10105e-16, 6.130983e-16, 
    6.123459e-16, 6.130629e-16, 6.128456e-16, 6.130657e-16, 6.119621e-16, 
    6.12435e-16, 6.114637e-16, 6.076747e-16, 6.087892e-16, 6.054625e-16, 
    6.03458e-16, 6.021265e-16, 6.011806e-16, 6.013143e-16, 6.015692e-16, 
    6.028788e-16, 6.041097e-16, 6.050469e-16, 6.056733e-16, 6.062905e-16, 
    6.081556e-16, 6.09143e-16, 6.113504e-16, 6.109526e-16, 6.116267e-16, 
    6.122711e-16, 6.133516e-16, 6.131739e-16, 6.136496e-16, 6.116093e-16, 
    6.129655e-16, 6.107263e-16, 6.113387e-16, 6.064564e-16, 6.045945e-16, 
    6.038009e-16, 6.031073e-16, 6.014171e-16, 6.025844e-16, 6.021243e-16, 
    6.03219e-16, 6.03914e-16, 6.035704e-16, 6.056905e-16, 6.048665e-16, 
    6.092015e-16, 6.073358e-16, 6.121959e-16, 6.110343e-16, 6.124743e-16, 
    6.117398e-16, 6.12998e-16, 6.118656e-16, 6.138268e-16, 6.142533e-16, 
    6.139619e-16, 6.150819e-16, 6.118028e-16, 6.130627e-16, 6.035607e-16, 
    6.036167e-16, 6.03878e-16, 6.027293e-16, 6.026591e-16, 6.016062e-16, 
    6.025432e-16, 6.029419e-16, 6.039544e-16, 6.045526e-16, 6.051212e-16, 
    6.063707e-16, 6.077645e-16, 6.097121e-16, 6.111097e-16, 6.120459e-16, 
    6.11472e-16, 6.119787e-16, 6.114122e-16, 6.111467e-16, 6.140934e-16, 
    6.124393e-16, 6.149208e-16, 6.147837e-16, 6.136609e-16, 6.147991e-16, 
    6.036561e-16, 6.033335e-16, 6.022127e-16, 6.030899e-16, 6.014915e-16, 
    6.023862e-16, 6.029003e-16, 6.048833e-16, 6.053191e-16, 6.057226e-16, 
    6.065195e-16, 6.075413e-16, 6.093322e-16, 6.108886e-16, 6.123086e-16, 
    6.122047e-16, 6.122412e-16, 6.125581e-16, 6.117728e-16, 6.12687e-16, 
    6.128402e-16, 6.124393e-16, 6.147653e-16, 6.141012e-16, 6.147807e-16, 
    6.143484e-16, 6.034384e-16, 6.039811e-16, 6.036879e-16, 6.042392e-16, 
    6.038507e-16, 6.055771e-16, 6.060943e-16, 6.085128e-16, 6.075211e-16, 
    6.090995e-16, 6.076817e-16, 6.079329e-16, 6.091501e-16, 6.077584e-16, 
    6.108024e-16, 6.087388e-16, 6.125704e-16, 6.105113e-16, 6.126994e-16, 
    6.123025e-16, 6.129597e-16, 6.135478e-16, 6.142878e-16, 6.156517e-16, 
    6.15336e-16, 6.164761e-16, 6.0479e-16, 6.054931e-16, 6.054316e-16, 
    6.061674e-16, 6.067112e-16, 6.078896e-16, 6.097774e-16, 6.090679e-16, 
    6.103706e-16, 6.106319e-16, 6.086529e-16, 6.09868e-16, 6.059638e-16, 
    6.065949e-16, 6.062195e-16, 6.048453e-16, 6.09231e-16, 6.069816e-16, 
    6.111327e-16, 6.099164e-16, 6.13464e-16, 6.117002e-16, 6.151621e-16, 
    6.166387e-16, 6.180287e-16, 6.196494e-16, 6.058772e-16, 6.053995e-16, 
    6.062549e-16, 6.07437e-16, 6.08534e-16, 6.099906e-16, 6.101397e-16, 
    6.104123e-16, 6.111183e-16, 6.117117e-16, 6.104982e-16, 6.118605e-16, 
    6.067406e-16, 6.094262e-16, 6.052185e-16, 6.064863e-16, 6.073675e-16, 
    6.069814e-16, 6.089869e-16, 6.094591e-16, 6.113759e-16, 6.103857e-16, 
    6.162741e-16, 6.136716e-16, 6.208835e-16, 6.188714e-16, 6.052325e-16, 
    6.058756e-16, 6.081114e-16, 6.070481e-16, 6.10088e-16, 6.108348e-16, 
    6.114423e-16, 6.122178e-16, 6.123018e-16, 6.127612e-16, 6.120083e-16, 
    6.127316e-16, 6.099937e-16, 6.112177e-16, 6.078565e-16, 6.086751e-16, 
    6.082987e-16, 6.078854e-16, 6.091605e-16, 6.105172e-16, 6.105467e-16, 
    6.109811e-16, 6.122043e-16, 6.101003e-16, 6.166086e-16, 6.125914e-16, 
    6.065767e-16, 6.078134e-16, 6.079906e-16, 6.075116e-16, 6.107603e-16, 
    6.095838e-16, 6.1275e-16, 6.11895e-16, 6.132958e-16, 6.125999e-16, 
    6.124974e-16, 6.116031e-16, 6.110459e-16, 6.096377e-16, 6.084909e-16, 
    6.075811e-16, 6.077928e-16, 6.08792e-16, 6.106003e-16, 6.123092e-16, 
    6.119348e-16, 6.131894e-16, 6.098677e-16, 6.11261e-16, 6.107227e-16, 
    6.121266e-16, 6.090489e-16, 6.116684e-16, 6.083784e-16, 6.086673e-16, 
    6.095605e-16, 6.113551e-16, 6.117527e-16, 6.121762e-16, 6.11915e-16, 
    6.106463e-16, 6.104385e-16, 6.095389e-16, 6.092902e-16, 6.086044e-16, 
    6.080362e-16, 6.085553e-16, 6.091e-16, 6.106471e-16, 6.120392e-16, 
    6.135562e-16, 6.139274e-16, 6.15696e-16, 6.142556e-16, 6.166309e-16, 
    6.146105e-16, 6.181067e-16, 6.118208e-16, 6.145522e-16, 6.096013e-16, 
    6.101356e-16, 6.111007e-16, 6.133137e-16, 6.1212e-16, 6.135162e-16, 
    6.104304e-16, 6.088261e-16, 6.084114e-16, 6.076363e-16, 6.084292e-16, 
    6.083647e-16, 6.09123e-16, 6.088794e-16, 6.106984e-16, 6.097216e-16, 
    6.124947e-16, 6.135053e-16, 6.163565e-16, 6.181012e-16, 6.198761e-16, 
    6.206586e-16, 6.208967e-16, 6.209962e-16 ;

 CWDC_TO_LITR2C =
  4.573201e-16, 4.585554e-16, 4.583154e-16, 4.593108e-16, 4.587589e-16, 
    4.594104e-16, 4.575709e-16, 4.586042e-16, 4.579448e-16, 4.574316e-16, 
    4.612395e-16, 4.593552e-16, 4.631953e-16, 4.619956e-16, 4.650072e-16, 
    4.630084e-16, 4.654099e-16, 4.649499e-16, 4.663347e-16, 4.659382e-16, 
    4.677066e-16, 4.665176e-16, 4.686229e-16, 4.67423e-16, 4.676106e-16, 
    4.664783e-16, 4.59735e-16, 4.61005e-16, 4.596597e-16, 4.598409e-16, 
    4.597597e-16, 4.587701e-16, 4.582709e-16, 4.572259e-16, 4.574158e-16, 
    4.581834e-16, 4.599224e-16, 4.593326e-16, 4.608192e-16, 4.607856e-16, 
    4.624381e-16, 4.616933e-16, 4.644673e-16, 4.636798e-16, 4.659547e-16, 
    4.653829e-16, 4.659278e-16, 4.657627e-16, 4.6593e-16, 4.650912e-16, 
    4.654506e-16, 4.647125e-16, 4.618328e-16, 4.626797e-16, 4.601515e-16, 
    4.586281e-16, 4.576161e-16, 4.568972e-16, 4.569989e-16, 4.571925e-16, 
    4.581879e-16, 4.591234e-16, 4.598356e-16, 4.603117e-16, 4.607808e-16, 
    4.621982e-16, 4.629487e-16, 4.646263e-16, 4.64324e-16, 4.648363e-16, 
    4.65326e-16, 4.661472e-16, 4.660122e-16, 4.663737e-16, 4.64823e-16, 
    4.658538e-16, 4.64152e-16, 4.646174e-16, 4.609069e-16, 4.594918e-16, 
    4.588887e-16, 4.583615e-16, 4.57077e-16, 4.579641e-16, 4.576145e-16, 
    4.584465e-16, 4.589746e-16, 4.587135e-16, 4.603248e-16, 4.596985e-16, 
    4.629931e-16, 4.615752e-16, 4.652689e-16, 4.643861e-16, 4.654804e-16, 
    4.649222e-16, 4.658784e-16, 4.650179e-16, 4.665084e-16, 4.668325e-16, 
    4.66611e-16, 4.674622e-16, 4.649702e-16, 4.659277e-16, 4.587061e-16, 
    4.587487e-16, 4.589472e-16, 4.580743e-16, 4.580209e-16, 4.572207e-16, 
    4.579329e-16, 4.582359e-16, 4.590054e-16, 4.5946e-16, 4.598921e-16, 
    4.608417e-16, 4.61901e-16, 4.633812e-16, 4.644433e-16, 4.651549e-16, 
    4.647187e-16, 4.651038e-16, 4.646733e-16, 4.644715e-16, 4.66711e-16, 
    4.654539e-16, 4.673398e-16, 4.672356e-16, 4.663823e-16, 4.672474e-16, 
    4.587786e-16, 4.585335e-16, 4.576816e-16, 4.583483e-16, 4.571335e-16, 
    4.578135e-16, 4.582042e-16, 4.597114e-16, 4.600425e-16, 4.603492e-16, 
    4.609548e-16, 4.617314e-16, 4.630924e-16, 4.642753e-16, 4.653546e-16, 
    4.652756e-16, 4.653034e-16, 4.655442e-16, 4.649473e-16, 4.656421e-16, 
    4.657585e-16, 4.654539e-16, 4.672216e-16, 4.667169e-16, 4.672334e-16, 
    4.669048e-16, 4.586132e-16, 4.590257e-16, 4.588028e-16, 4.592218e-16, 
    4.589265e-16, 4.602386e-16, 4.606317e-16, 4.624697e-16, 4.617161e-16, 
    4.629156e-16, 4.61838e-16, 4.62029e-16, 4.629541e-16, 4.618964e-16, 
    4.642099e-16, 4.626415e-16, 4.655536e-16, 4.639886e-16, 4.656515e-16, 
    4.653499e-16, 4.658494e-16, 4.662964e-16, 4.668587e-16, 4.678952e-16, 
    4.676554e-16, 4.685219e-16, 4.596404e-16, 4.601748e-16, 4.60128e-16, 
    4.606872e-16, 4.611005e-16, 4.619961e-16, 4.634309e-16, 4.628916e-16, 
    4.638817e-16, 4.640802e-16, 4.625762e-16, 4.634997e-16, 4.605325e-16, 
    4.610121e-16, 4.607268e-16, 4.596825e-16, 4.630156e-16, 4.61306e-16, 
    4.644608e-16, 4.635365e-16, 4.662326e-16, 4.648922e-16, 4.675232e-16, 
    4.686454e-16, 4.697018e-16, 4.709336e-16, 4.604666e-16, 4.601036e-16, 
    4.607537e-16, 4.616521e-16, 4.624858e-16, 4.635929e-16, 4.637062e-16, 
    4.639134e-16, 4.644499e-16, 4.649009e-16, 4.639786e-16, 4.65014e-16, 
    4.611228e-16, 4.63164e-16, 4.599661e-16, 4.609297e-16, 4.615993e-16, 
    4.613058e-16, 4.6283e-16, 4.631889e-16, 4.646457e-16, 4.638931e-16, 
    4.683684e-16, 4.663904e-16, 4.718714e-16, 4.703423e-16, 4.599767e-16, 
    4.604655e-16, 4.621647e-16, 4.613566e-16, 4.636668e-16, 4.642345e-16, 
    4.646961e-16, 4.652855e-16, 4.653494e-16, 4.656984e-16, 4.651263e-16, 
    4.65676e-16, 4.635952e-16, 4.645254e-16, 4.619709e-16, 4.625931e-16, 
    4.62307e-16, 4.619929e-16, 4.62962e-16, 4.639931e-16, 4.640156e-16, 
    4.643456e-16, 4.652753e-16, 4.636762e-16, 4.686226e-16, 4.655694e-16, 
    4.609983e-16, 4.619382e-16, 4.620728e-16, 4.617088e-16, 4.641778e-16, 
    4.632837e-16, 4.6569e-16, 4.650402e-16, 4.661048e-16, 4.655759e-16, 
    4.65498e-16, 4.648183e-16, 4.643949e-16, 4.633246e-16, 4.62453e-16, 
    4.617617e-16, 4.619225e-16, 4.626818e-16, 4.640562e-16, 4.653549e-16, 
    4.650705e-16, 4.66024e-16, 4.634995e-16, 4.645583e-16, 4.641492e-16, 
    4.652162e-16, 4.628772e-16, 4.648679e-16, 4.623676e-16, 4.625871e-16, 
    4.63266e-16, 4.646299e-16, 4.649321e-16, 4.652539e-16, 4.650554e-16, 
    4.640912e-16, 4.639333e-16, 4.632496e-16, 4.630605e-16, 4.625394e-16, 
    4.621075e-16, 4.62502e-16, 4.62916e-16, 4.640918e-16, 4.651498e-16, 
    4.663027e-16, 4.665848e-16, 4.679289e-16, 4.668343e-16, 4.686395e-16, 
    4.67104e-16, 4.697611e-16, 4.649838e-16, 4.670597e-16, 4.63297e-16, 
    4.637031e-16, 4.644365e-16, 4.661184e-16, 4.652111e-16, 4.662723e-16, 
    4.639271e-16, 4.627078e-16, 4.623927e-16, 4.618036e-16, 4.624062e-16, 
    4.623572e-16, 4.629335e-16, 4.627483e-16, 4.641308e-16, 4.633884e-16, 
    4.65496e-16, 4.662641e-16, 4.684309e-16, 4.69757e-16, 4.711058e-16, 
    4.717005e-16, 4.718815e-16, 4.719571e-16 ;

 CWDC_TO_LITR3C =
  1.444169e-16, 1.44807e-16, 1.447312e-16, 1.450455e-16, 1.448712e-16, 
    1.45077e-16, 1.444961e-16, 1.448224e-16, 1.446141e-16, 1.444521e-16, 
    1.456546e-16, 1.450595e-16, 1.462722e-16, 1.458934e-16, 1.468444e-16, 
    1.462132e-16, 1.469715e-16, 1.468263e-16, 1.472636e-16, 1.471384e-16, 
    1.476968e-16, 1.473214e-16, 1.479862e-16, 1.476073e-16, 1.476665e-16, 
    1.473089e-16, 1.451795e-16, 1.455805e-16, 1.451557e-16, 1.452129e-16, 
    1.451873e-16, 1.448748e-16, 1.447171e-16, 1.443871e-16, 1.444471e-16, 
    1.446895e-16, 1.452386e-16, 1.450524e-16, 1.455218e-16, 1.455112e-16, 
    1.460331e-16, 1.457979e-16, 1.466739e-16, 1.464252e-16, 1.471436e-16, 
    1.46963e-16, 1.471351e-16, 1.470829e-16, 1.471358e-16, 1.468709e-16, 
    1.469844e-16, 1.467513e-16, 1.458419e-16, 1.461094e-16, 1.45311e-16, 
    1.448299e-16, 1.445104e-16, 1.442833e-16, 1.443154e-16, 1.443766e-16, 
    1.446909e-16, 1.449863e-16, 1.452112e-16, 1.453616e-16, 1.455097e-16, 
    1.459573e-16, 1.461943e-16, 1.467241e-16, 1.466286e-16, 1.467904e-16, 
    1.469451e-16, 1.472044e-16, 1.471617e-16, 1.472759e-16, 1.467862e-16, 
    1.471117e-16, 1.465743e-16, 1.467213e-16, 1.455495e-16, 1.451027e-16, 
    1.449122e-16, 1.447457e-16, 1.443401e-16, 1.446202e-16, 1.445098e-16, 
    1.447726e-16, 1.449394e-16, 1.448569e-16, 1.453657e-16, 1.45168e-16, 
    1.462084e-16, 1.457606e-16, 1.46927e-16, 1.466482e-16, 1.469938e-16, 
    1.468175e-16, 1.471195e-16, 1.468478e-16, 1.473184e-16, 1.474208e-16, 
    1.473508e-16, 1.476196e-16, 1.468327e-16, 1.47135e-16, 1.448546e-16, 
    1.44868e-16, 1.449307e-16, 1.44655e-16, 1.446382e-16, 1.443855e-16, 
    1.446104e-16, 1.447061e-16, 1.449491e-16, 1.450926e-16, 1.452291e-16, 
    1.45529e-16, 1.458635e-16, 1.463309e-16, 1.466663e-16, 1.46891e-16, 
    1.467533e-16, 1.468749e-16, 1.467389e-16, 1.466752e-16, 1.473824e-16, 
    1.469854e-16, 1.47581e-16, 1.475481e-16, 1.472786e-16, 1.475518e-16, 
    1.448775e-16, 1.448001e-16, 1.44531e-16, 1.447416e-16, 1.44358e-16, 
    1.445727e-16, 1.446961e-16, 1.45172e-16, 1.452766e-16, 1.453734e-16, 
    1.455647e-16, 1.458099e-16, 1.462397e-16, 1.466133e-16, 1.469541e-16, 
    1.469291e-16, 1.469379e-16, 1.47014e-16, 1.468255e-16, 1.470449e-16, 
    1.470816e-16, 1.469854e-16, 1.475437e-16, 1.473843e-16, 1.475474e-16, 
    1.474436e-16, 1.448252e-16, 1.449555e-16, 1.448851e-16, 1.450174e-16, 
    1.449242e-16, 1.453385e-16, 1.454626e-16, 1.460431e-16, 1.458051e-16, 
    1.461839e-16, 1.458436e-16, 1.459039e-16, 1.46196e-16, 1.45862e-16, 
    1.465926e-16, 1.460973e-16, 1.470169e-16, 1.465227e-16, 1.470478e-16, 
    1.469526e-16, 1.471103e-16, 1.472515e-16, 1.474291e-16, 1.477564e-16, 
    1.476806e-16, 1.479543e-16, 1.451496e-16, 1.453184e-16, 1.453036e-16, 
    1.454802e-16, 1.456107e-16, 1.458935e-16, 1.463466e-16, 1.461763e-16, 
    1.464889e-16, 1.465517e-16, 1.460767e-16, 1.463683e-16, 1.454313e-16, 
    1.455828e-16, 1.454927e-16, 1.451629e-16, 1.462154e-16, 1.456756e-16, 
    1.466718e-16, 1.463799e-16, 1.472314e-16, 1.468081e-16, 1.476389e-16, 
    1.479933e-16, 1.483269e-16, 1.487159e-16, 1.454105e-16, 1.452959e-16, 
    1.455012e-16, 1.457849e-16, 1.460482e-16, 1.463977e-16, 1.464335e-16, 
    1.46499e-16, 1.466684e-16, 1.468108e-16, 1.465196e-16, 1.468465e-16, 
    1.456177e-16, 1.462623e-16, 1.452525e-16, 1.455567e-16, 1.457682e-16, 
    1.456755e-16, 1.461569e-16, 1.462702e-16, 1.467302e-16, 1.464926e-16, 
    1.479058e-16, 1.472812e-16, 1.49012e-16, 1.485291e-16, 1.452558e-16, 
    1.454102e-16, 1.459467e-16, 1.456915e-16, 1.464211e-16, 1.466004e-16, 
    1.467461e-16, 1.469323e-16, 1.469524e-16, 1.470627e-16, 1.46882e-16, 
    1.470556e-16, 1.463985e-16, 1.466922e-16, 1.458855e-16, 1.46082e-16, 
    1.459917e-16, 1.458925e-16, 1.461985e-16, 1.465241e-16, 1.465312e-16, 
    1.466355e-16, 1.46929e-16, 1.464241e-16, 1.479861e-16, 1.470219e-16, 
    1.455784e-16, 1.458752e-16, 1.459177e-16, 1.458028e-16, 1.465825e-16, 
    1.463001e-16, 1.4706e-16, 1.468548e-16, 1.47191e-16, 1.47024e-16, 
    1.469994e-16, 1.467847e-16, 1.46651e-16, 1.46313e-16, 1.460378e-16, 
    1.458195e-16, 1.458703e-16, 1.461101e-16, 1.465441e-16, 1.469542e-16, 
    1.468644e-16, 1.471655e-16, 1.463683e-16, 1.467026e-16, 1.465734e-16, 
    1.469104e-16, 1.461717e-16, 1.468004e-16, 1.460108e-16, 1.460801e-16, 
    1.462945e-16, 1.467252e-16, 1.468207e-16, 1.469223e-16, 1.468596e-16, 
    1.465551e-16, 1.465052e-16, 1.462893e-16, 1.462297e-16, 1.460651e-16, 
    1.459287e-16, 1.460533e-16, 1.46184e-16, 1.465553e-16, 1.468894e-16, 
    1.472535e-16, 1.473426e-16, 1.47767e-16, 1.474213e-16, 1.479914e-16, 
    1.475065e-16, 1.483456e-16, 1.46837e-16, 1.474925e-16, 1.463043e-16, 
    1.464326e-16, 1.466642e-16, 1.471953e-16, 1.469088e-16, 1.472439e-16, 
    1.465033e-16, 1.461183e-16, 1.460188e-16, 1.458327e-16, 1.46023e-16, 
    1.460075e-16, 1.461895e-16, 1.461311e-16, 1.465676e-16, 1.463332e-16, 
    1.469987e-16, 1.472413e-16, 1.479256e-16, 1.483443e-16, 1.487702e-16, 
    1.489581e-16, 1.490152e-16, 1.490391e-16 ;

 CWDC_vr =
  5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110344e-05, 5.110345e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110345e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 
    5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 
    5.110343e-05, 5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110345e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110343e-05, 5.110344e-05, 5.110343e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110342e-05, 5.110343e-05, 5.110343e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 5.110344e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDN =
  1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.78993e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789931e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09 ;

 CWDN_TO_LITR2N =
  9.146403e-19, 9.171108e-19, 9.166309e-19, 9.186216e-19, 9.175177e-19, 
    9.188207e-19, 9.151418e-19, 9.172085e-19, 9.158895e-19, 9.148633e-19, 
    9.224791e-19, 9.187104e-19, 9.263906e-19, 9.239912e-19, 9.300143e-19, 
    9.260169e-19, 9.308197e-19, 9.298999e-19, 9.326693e-19, 9.318763e-19, 
    9.354132e-19, 9.330352e-19, 9.372458e-19, 9.348459e-19, 9.352213e-19, 
    9.329566e-19, 9.194701e-19, 9.220099e-19, 9.193193e-19, 9.196817e-19, 
    9.195193e-19, 9.175403e-19, 9.165419e-19, 9.144519e-19, 9.148317e-19, 
    9.163669e-19, 9.198447e-19, 9.186652e-19, 9.216383e-19, 9.215712e-19, 
    9.248761e-19, 9.233866e-19, 9.289346e-19, 9.273596e-19, 9.319094e-19, 
    9.307658e-19, 9.318556e-19, 9.315253e-19, 9.318599e-19, 9.301824e-19, 
    9.309012e-19, 9.294249e-19, 9.236654e-19, 9.253595e-19, 9.203031e-19, 
    9.172561e-19, 9.152322e-19, 9.137945e-19, 9.139978e-19, 9.143851e-19, 
    9.163758e-19, 9.182467e-19, 9.196712e-19, 9.206235e-19, 9.215615e-19, 
    9.243965e-19, 9.258974e-19, 9.292526e-19, 9.286481e-19, 9.296726e-19, 
    9.30652e-19, 9.322945e-19, 9.320243e-19, 9.327475e-19, 9.296461e-19, 
    9.317075e-19, 9.28304e-19, 9.292348e-19, 9.218138e-19, 9.189836e-19, 
    9.177774e-19, 9.16723e-19, 9.14154e-19, 9.159283e-19, 9.152289e-19, 
    9.168929e-19, 9.179492e-19, 9.174269e-19, 9.206495e-19, 9.193971e-19, 
    9.259863e-19, 9.231504e-19, 9.305379e-19, 9.287721e-19, 9.30961e-19, 
    9.298445e-19, 9.317569e-19, 9.300358e-19, 9.330168e-19, 9.33665e-19, 
    9.332221e-19, 9.349244e-19, 9.299402e-19, 9.318554e-19, 9.174122e-19, 
    9.174974e-19, 9.178945e-19, 9.161484e-19, 9.160417e-19, 9.144413e-19, 
    9.158657e-19, 9.164718e-19, 9.180107e-19, 9.1892e-19, 9.197842e-19, 
    9.216834e-19, 9.23802e-19, 9.267623e-19, 9.288866e-19, 9.303098e-19, 
    9.294374e-19, 9.302076e-19, 9.293465e-19, 9.28943e-19, 9.33422e-19, 
    9.309077e-19, 9.346797e-19, 9.344712e-19, 9.327645e-19, 9.344947e-19, 
    9.175572e-19, 9.17067e-19, 9.153632e-19, 9.166967e-19, 9.14267e-19, 
    9.15627e-19, 9.164084e-19, 9.194227e-19, 9.200851e-19, 9.206983e-19, 
    9.219096e-19, 9.234628e-19, 9.261849e-19, 9.285507e-19, 9.307091e-19, 
    9.305511e-19, 9.306067e-19, 9.310884e-19, 9.298947e-19, 9.312843e-19, 
    9.315171e-19, 9.309078e-19, 9.344432e-19, 9.334338e-19, 9.344668e-19, 
    9.338096e-19, 9.172265e-19, 9.180514e-19, 9.176056e-19, 9.184436e-19, 
    9.17853e-19, 9.204772e-19, 9.212633e-19, 9.249394e-19, 9.234321e-19, 
    9.258312e-19, 9.236761e-19, 9.240579e-19, 9.259082e-19, 9.237928e-19, 
    9.284198e-19, 9.25283e-19, 9.311071e-19, 9.279771e-19, 9.31303e-19, 
    9.306998e-19, 9.316987e-19, 9.325928e-19, 9.337174e-19, 9.357905e-19, 
    9.353107e-19, 9.370437e-19, 9.192809e-19, 9.203496e-19, 9.20256e-19, 
    9.213744e-19, 9.22201e-19, 9.239923e-19, 9.268618e-19, 9.257832e-19, 
    9.277634e-19, 9.281604e-19, 9.251524e-19, 9.269993e-19, 9.21065e-19, 
    9.220242e-19, 9.214536e-19, 9.193648e-19, 9.260311e-19, 9.22612e-19, 
    9.289217e-19, 9.27073e-19, 9.324652e-19, 9.297843e-19, 9.350465e-19, 
    9.372909e-19, 9.394036e-19, 9.418671e-19, 9.209333e-19, 9.202072e-19, 
    9.215075e-19, 9.233043e-19, 9.249717e-19, 9.271857e-19, 9.274125e-19, 
    9.278268e-19, 9.288998e-19, 9.298019e-19, 9.279573e-19, 9.30028e-19, 
    9.222456e-19, 9.263279e-19, 9.199322e-19, 9.218593e-19, 9.231986e-19, 
    9.226117e-19, 9.256601e-19, 9.263778e-19, 9.292913e-19, 9.277862e-19, 
    9.367367e-19, 9.327808e-19, 9.437429e-19, 9.406846e-19, 9.199534e-19, 
    9.20931e-19, 9.243294e-19, 9.227131e-19, 9.273337e-19, 9.284689e-19, 
    9.293922e-19, 9.305711e-19, 9.306988e-19, 9.313969e-19, 9.302526e-19, 
    9.313519e-19, 9.271905e-19, 9.290508e-19, 9.239418e-19, 9.251862e-19, 
    9.24614e-19, 9.239858e-19, 9.25924e-19, 9.279862e-19, 9.280311e-19, 
    9.286913e-19, 9.305506e-19, 9.273524e-19, 9.372452e-19, 9.311389e-19, 
    9.219965e-19, 9.238764e-19, 9.241457e-19, 9.234176e-19, 9.283556e-19, 
    9.265675e-19, 9.3138e-19, 9.300804e-19, 9.322097e-19, 9.311517e-19, 
    9.30996e-19, 9.296368e-19, 9.287898e-19, 9.266493e-19, 9.249061e-19, 
    9.235233e-19, 9.238449e-19, 9.253637e-19, 9.281125e-19, 9.307099e-19, 
    9.301409e-19, 9.320479e-19, 9.26999e-19, 9.291167e-19, 9.282985e-19, 
    9.304324e-19, 9.257544e-19, 9.297359e-19, 9.247352e-19, 9.251742e-19, 
    9.265319e-19, 9.292598e-19, 9.298641e-19, 9.305079e-19, 9.301108e-19, 
    9.281824e-19, 9.278666e-19, 9.264992e-19, 9.261211e-19, 9.250788e-19, 
    9.24215e-19, 9.250039e-19, 9.25832e-19, 9.281835e-19, 9.302996e-19, 
    9.326054e-19, 9.331695e-19, 9.358579e-19, 9.336685e-19, 9.37279e-19, 
    9.34208e-19, 9.395222e-19, 9.299676e-19, 9.341193e-19, 9.26594e-19, 
    9.274062e-19, 9.288731e-19, 9.322368e-19, 9.304224e-19, 9.325446e-19, 
    9.278543e-19, 9.254157e-19, 9.247854e-19, 9.236072e-19, 9.248123e-19, 
    9.247144e-19, 9.25867e-19, 9.254967e-19, 9.282616e-19, 9.267768e-19, 
    9.309919e-19, 9.325281e-19, 9.368619e-19, 9.395139e-19, 9.422116e-19, 
    9.43401e-19, 9.43763e-19, 9.439143e-19 ;

 CWDN_TO_LITR3N =
  2.888338e-19, 2.896139e-19, 2.894624e-19, 2.90091e-19, 2.897424e-19, 
    2.901539e-19, 2.889921e-19, 2.896448e-19, 2.892283e-19, 2.889042e-19, 
    2.913092e-19, 2.901191e-19, 2.925444e-19, 2.917867e-19, 2.936887e-19, 
    2.924264e-19, 2.939431e-19, 2.936526e-19, 2.945271e-19, 2.942767e-19, 
    2.953936e-19, 2.946427e-19, 2.959723e-19, 2.952145e-19, 2.95333e-19, 
    2.946179e-19, 2.90359e-19, 2.91161e-19, 2.903114e-19, 2.904258e-19, 
    2.903745e-19, 2.897496e-19, 2.894343e-19, 2.887743e-19, 2.888942e-19, 
    2.89379e-19, 2.904773e-19, 2.901048e-19, 2.910437e-19, 2.910225e-19, 
    2.920662e-19, 2.915957e-19, 2.933477e-19, 2.928504e-19, 2.942872e-19, 
    2.93926e-19, 2.942702e-19, 2.941659e-19, 2.942715e-19, 2.937418e-19, 
    2.939688e-19, 2.935026e-19, 2.916838e-19, 2.922188e-19, 2.90622e-19, 
    2.896598e-19, 2.890207e-19, 2.885667e-19, 2.886309e-19, 2.887532e-19, 
    2.893818e-19, 2.899726e-19, 2.904225e-19, 2.907232e-19, 2.910194e-19, 
    2.919147e-19, 2.923886e-19, 2.934482e-19, 2.932573e-19, 2.935808e-19, 
    2.938901e-19, 2.944088e-19, 2.943235e-19, 2.945518e-19, 2.935724e-19, 
    2.942234e-19, 2.931486e-19, 2.934426e-19, 2.910991e-19, 2.902054e-19, 
    2.898244e-19, 2.894915e-19, 2.886802e-19, 2.892405e-19, 2.890197e-19, 
    2.895451e-19, 2.898787e-19, 2.897138e-19, 2.907314e-19, 2.903359e-19, 
    2.924167e-19, 2.915212e-19, 2.938541e-19, 2.932965e-19, 2.939877e-19, 
    2.936351e-19, 2.94239e-19, 2.936955e-19, 2.946369e-19, 2.948416e-19, 
    2.947017e-19, 2.952393e-19, 2.936654e-19, 2.942701e-19, 2.897091e-19, 
    2.89736e-19, 2.898614e-19, 2.8931e-19, 2.892764e-19, 2.887709e-19, 
    2.892208e-19, 2.894121e-19, 2.898981e-19, 2.901852e-19, 2.904582e-19, 
    2.910579e-19, 2.91727e-19, 2.926618e-19, 2.933326e-19, 2.93782e-19, 
    2.935066e-19, 2.937497e-19, 2.934778e-19, 2.933504e-19, 2.947649e-19, 
    2.939709e-19, 2.95162e-19, 2.950962e-19, 2.945572e-19, 2.951036e-19, 
    2.897549e-19, 2.896001e-19, 2.890621e-19, 2.894832e-19, 2.887159e-19, 
    2.891454e-19, 2.893921e-19, 2.90344e-19, 2.905532e-19, 2.907469e-19, 
    2.911293e-19, 2.916198e-19, 2.924794e-19, 2.932265e-19, 2.939082e-19, 
    2.938582e-19, 2.938758e-19, 2.940279e-19, 2.93651e-19, 2.940898e-19, 
    2.941633e-19, 2.939709e-19, 2.950873e-19, 2.947686e-19, 2.950948e-19, 
    2.948873e-19, 2.896504e-19, 2.89911e-19, 2.897702e-19, 2.900348e-19, 
    2.898483e-19, 2.90677e-19, 2.909253e-19, 2.920861e-19, 2.916101e-19, 
    2.923678e-19, 2.916872e-19, 2.918078e-19, 2.923921e-19, 2.91724e-19, 
    2.931852e-19, 2.921946e-19, 2.940338e-19, 2.930454e-19, 2.940957e-19, 
    2.939052e-19, 2.942206e-19, 2.94503e-19, 2.948581e-19, 2.955128e-19, 
    2.953613e-19, 2.959085e-19, 2.902992e-19, 2.906367e-19, 2.906072e-19, 
    2.909603e-19, 2.912214e-19, 2.91787e-19, 2.926932e-19, 2.923526e-19, 
    2.929779e-19, 2.931033e-19, 2.921534e-19, 2.927366e-19, 2.908626e-19, 
    2.911656e-19, 2.909853e-19, 2.903257e-19, 2.924309e-19, 2.913512e-19, 
    2.933437e-19, 2.927599e-19, 2.944627e-19, 2.936161e-19, 2.952778e-19, 
    2.959866e-19, 2.966538e-19, 2.974317e-19, 2.90821e-19, 2.905918e-19, 
    2.910024e-19, 2.915698e-19, 2.920963e-19, 2.927955e-19, 2.928671e-19, 
    2.929979e-19, 2.933368e-19, 2.936216e-19, 2.930391e-19, 2.93693e-19, 
    2.912355e-19, 2.925246e-19, 2.905049e-19, 2.911134e-19, 2.915364e-19, 
    2.913511e-19, 2.923137e-19, 2.925404e-19, 2.934604e-19, 2.929851e-19, 
    2.958116e-19, 2.945624e-19, 2.98024e-19, 2.970583e-19, 2.905116e-19, 
    2.908203e-19, 2.918935e-19, 2.913831e-19, 2.928422e-19, 2.932007e-19, 
    2.934923e-19, 2.938645e-19, 2.939048e-19, 2.941253e-19, 2.93764e-19, 
    2.941111e-19, 2.92797e-19, 2.933845e-19, 2.917711e-19, 2.92164e-19, 
    2.919834e-19, 2.91785e-19, 2.92397e-19, 2.930483e-19, 2.930624e-19, 
    2.932709e-19, 2.938581e-19, 2.928481e-19, 2.959722e-19, 2.940439e-19, 
    2.911568e-19, 2.917504e-19, 2.918355e-19, 2.916056e-19, 2.931649e-19, 
    2.926003e-19, 2.9412e-19, 2.937096e-19, 2.94382e-19, 2.940479e-19, 
    2.939988e-19, 2.935695e-19, 2.93302e-19, 2.926261e-19, 2.920756e-19, 
    2.916389e-19, 2.917405e-19, 2.922201e-19, 2.930881e-19, 2.939084e-19, 
    2.937287e-19, 2.943309e-19, 2.927365e-19, 2.934053e-19, 2.931469e-19, 
    2.938207e-19, 2.923435e-19, 2.936008e-19, 2.920216e-19, 2.921603e-19, 
    2.92589e-19, 2.934504e-19, 2.936413e-19, 2.938446e-19, 2.937192e-19, 
    2.931102e-19, 2.930105e-19, 2.925787e-19, 2.924593e-19, 2.921301e-19, 
    2.918574e-19, 2.921065e-19, 2.92368e-19, 2.931106e-19, 2.937788e-19, 
    2.94507e-19, 2.946851e-19, 2.955341e-19, 2.948427e-19, 2.959828e-19, 
    2.950131e-19, 2.966912e-19, 2.93674e-19, 2.949851e-19, 2.926086e-19, 
    2.928651e-19, 2.933283e-19, 2.943906e-19, 2.938176e-19, 2.944878e-19, 
    2.930066e-19, 2.922365e-19, 2.920375e-19, 2.916655e-19, 2.92046e-19, 
    2.920151e-19, 2.92379e-19, 2.922621e-19, 2.931352e-19, 2.926664e-19, 
    2.939974e-19, 2.944826e-19, 2.958511e-19, 2.966886e-19, 2.975405e-19, 
    2.979161e-19, 2.980304e-19, 2.980782e-19 ;

 CWDN_vr =
  1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADSTEMC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 DEADSTEMN =
  6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05 ;

 DENIT =
  2.809608e-14, 2.822132e-14, 2.81969e-14, 2.8298e-14, 2.824186e-14, 
    2.830805e-14, 2.812131e-14, 2.822615e-14, 2.815916e-14, 2.81071e-14, 
    2.849427e-14, 2.830232e-14, 2.869362e-14, 2.857102e-14, 2.887894e-14, 
    2.867451e-14, 2.892015e-14, 2.887291e-14, 2.901485e-14, 2.897413e-14, 
    2.91559e-14, 2.903356e-14, 2.925006e-14, 2.91266e-14, 2.91459e-14, 
    2.902941e-14, 2.834104e-14, 2.847056e-14, 2.833334e-14, 2.83518e-14, 
    2.834347e-14, 2.824293e-14, 2.819234e-14, 2.808624e-14, 2.810545e-14, 
    2.818333e-14, 2.835992e-14, 2.829987e-14, 2.845101e-14, 2.84476e-14, 
    2.861606e-14, 2.854006e-14, 2.882346e-14, 2.874281e-14, 2.89758e-14, 
    2.891714e-14, 2.897301e-14, 2.895601e-14, 2.897315e-14, 2.88872e-14, 
    2.892397e-14, 2.884833e-14, 2.85546e-14, 2.864101e-14, 2.838332e-14, 
    2.822863e-14, 2.812581e-14, 2.805297e-14, 2.806321e-14, 2.808286e-14, 
    2.818374e-14, 2.827859e-14, 2.835094e-14, 2.839934e-14, 2.844704e-14, 
    2.859176e-14, 2.866824e-14, 2.883974e-14, 2.880871e-14, 2.886118e-14, 
    2.891128e-14, 2.899547e-14, 2.898159e-14, 2.901868e-14, 2.885963e-14, 
    2.896532e-14, 2.879083e-14, 2.883854e-14, 2.846047e-14, 2.831616e-14, 
    2.825504e-14, 2.820137e-14, 2.807112e-14, 2.816105e-14, 2.812557e-14, 
    2.820984e-14, 2.826346e-14, 2.823689e-14, 2.840064e-14, 2.833692e-14, 
    2.867274e-14, 2.8528e-14, 2.890547e-14, 2.881501e-14, 2.892707e-14, 
    2.886986e-14, 2.896786e-14, 2.887962e-14, 2.903243e-14, 2.906577e-14, 
    2.904294e-14, 2.913036e-14, 2.887457e-14, 2.897278e-14, 2.82363e-14, 
    2.824063e-14, 2.826075e-14, 2.817219e-14, 2.816675e-14, 2.808558e-14, 
    2.815772e-14, 2.818848e-14, 2.826649e-14, 2.831267e-14, 2.835656e-14, 
    2.84532e-14, 2.856119e-14, 2.871226e-14, 2.882085e-14, 2.889366e-14, 
    2.884896e-14, 2.888837e-14, 2.884427e-14, 2.882356e-14, 2.905322e-14, 
    2.892423e-14, 2.911771e-14, 2.9107e-14, 2.901938e-14, 2.910813e-14, 
    2.824362e-14, 2.821868e-14, 2.813231e-14, 2.819985e-14, 2.807669e-14, 
    2.814563e-14, 2.818527e-14, 2.833826e-14, 2.837182e-14, 2.840305e-14, 
    2.846465e-14, 2.854377e-14, 2.868271e-14, 2.880364e-14, 2.891409e-14, 
    2.890595e-14, 2.890879e-14, 2.893346e-14, 2.887228e-14, 2.894345e-14, 
    2.895539e-14, 2.892413e-14, 2.910549e-14, 2.905365e-14, 2.910667e-14, 
    2.907286e-14, 2.822674e-14, 2.82686e-14, 2.824593e-14, 2.828852e-14, 
    2.825848e-14, 2.839191e-14, 2.84319e-14, 2.861922e-14, 2.854222e-14, 
    2.866468e-14, 2.855459e-14, 2.85741e-14, 2.866868e-14, 2.856045e-14, 
    2.879692e-14, 2.86366e-14, 2.893439e-14, 2.877425e-14, 2.894438e-14, 
    2.891341e-14, 2.896458e-14, 2.901049e-14, 2.906815e-14, 2.917476e-14, 
    2.915e-14, 2.923916e-14, 2.833103e-14, 2.838539e-14, 2.838055e-14, 
    2.843742e-14, 2.847951e-14, 2.857078e-14, 2.871728e-14, 2.866211e-14, 
    2.876326e-14, 2.87836e-14, 2.862981e-14, 2.872423e-14, 2.842152e-14, 
    2.847038e-14, 2.844123e-14, 2.833496e-14, 2.867466e-14, 2.850022e-14, 
    2.882235e-14, 2.872773e-14, 2.900387e-14, 2.886652e-14, 2.91364e-14, 
    2.925202e-14, 2.936066e-14, 2.948791e-14, 2.841501e-14, 2.837801e-14, 
    2.844413e-14, 2.853579e-14, 2.86207e-14, 2.87338e-14, 2.874532e-14, 
    2.876649e-14, 2.882135e-14, 2.886755e-14, 2.877317e-14, 2.887905e-14, 
    2.848178e-14, 2.868978e-14, 2.836375e-14, 2.84619e-14, 2.853002e-14, 
    2.850008e-14, 2.865548e-14, 2.869211e-14, 2.884117e-14, 2.876407e-14, 
    2.922344e-14, 2.902005e-14, 2.95847e-14, 2.942677e-14, 2.836508e-14, 
    2.841476e-14, 2.858796e-14, 2.850551e-14, 2.874126e-14, 2.879937e-14, 
    2.884654e-14, 2.890698e-14, 2.891343e-14, 2.894924e-14, 2.889051e-14, 
    2.894686e-14, 2.873377e-14, 2.882894e-14, 2.856783e-14, 2.863132e-14, 
    2.860207e-14, 2.856999e-14, 2.866887e-14, 2.877439e-14, 2.877655e-14, 
    2.881037e-14, 2.890591e-14, 2.874176e-14, 2.924972e-14, 2.893592e-14, 
    2.846897e-14, 2.856487e-14, 2.857847e-14, 2.854132e-14, 2.879348e-14, 
    2.870206e-14, 2.894836e-14, 2.88817e-14, 2.899082e-14, 2.893659e-14, 
    2.892856e-14, 2.885891e-14, 2.881552e-14, 2.870607e-14, 2.861699e-14, 
    2.854641e-14, 2.856276e-14, 2.864032e-14, 2.878076e-14, 2.891373e-14, 
    2.888458e-14, 2.898221e-14, 2.872365e-14, 2.883205e-14, 2.879011e-14, 
    2.889933e-14, 2.866056e-14, 2.886451e-14, 2.860846e-14, 2.863084e-14, 
    2.870018e-14, 2.883982e-14, 2.887058e-14, 2.890361e-14, 2.888316e-14, 
    2.87845e-14, 2.876828e-14, 2.869831e-14, 2.867901e-14, 2.862573e-14, 
    2.858161e-14, 2.862189e-14, 2.866416e-14, 2.878432e-14, 2.889267e-14, 
    2.901084e-14, 2.903975e-14, 2.91781e-14, 2.906551e-14, 2.925136e-14, 
    2.909343e-14, 2.936677e-14, 2.887617e-14, 2.908917e-14, 2.870332e-14, 
    2.874479e-14, 2.881995e-14, 2.899231e-14, 2.889912e-14, 2.900805e-14, 
    2.876762e-14, 2.864306e-14, 2.861075e-14, 2.855067e-14, 2.861208e-14, 
    2.860708e-14, 2.866588e-14, 2.864693e-14, 2.878824e-14, 2.87123e-14, 
    2.892804e-14, 2.900687e-14, 2.922955e-14, 2.936619e-14, 2.95053e-14, 
    2.956674e-14, 2.958544e-14, 2.959324e-14 ;

 DISPVEGC =
  0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653 ;

 DISPVEGN =
  0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997 ;

 DSTDEP =
  2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12 ;

 DSTFLXT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_NFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_GRND_LAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 EFLX_LH_TOT =
  5.945704, 5.96459, 5.960935, 5.976095, 5.967731, 5.977613, 5.949567, 
    5.965309, 5.955278, 5.947451, 6.005329, 5.976777, 6.035303, 6.017036, 
    6.064812, 6.032414, 6.071017, 6.064003, 6.08531, 6.079208, 6.106329, 
    6.088128, 6.12053, 6.102022, 6.104887, 6.087515, 5.982594, 6.001753, 
    5.981442, 5.984177, 5.982967, 5.967877, 5.960184, 5.944315, 5.947209, 
    5.958894, 5.985409, 5.976478, 5.999142, 5.998631, 6.023797, 6.012445, 
    6.056595, 6.0428, 6.079464, 6.070662, 6.079037, 6.076507, 6.079071, 
    6.066167, 6.07169, 6.060366, 6.014556, 6.027471, 5.988921, 5.965604, 
    5.950243, 5.939291, 5.940838, 5.943774, 5.958961, 5.973293, 5.984146, 
    5.991398, 5.998557, 6.020007, 6.031534, 6.058997, 6.054414, 6.062228, 
    6.069789, 6.082406, 6.080338, 6.085884, 6.062068, 6.077869, 6.050041, 
    6.058909, 6.000245, 5.978899, 5.969609, 5.961628, 5.942023, 5.955546, 
    5.950208, 5.962965, 5.971028, 5.967055, 5.991597, 5.982049, 6.032218, 
    6.010608, 6.068908, 6.05536, 6.072166, 6.0636, 6.07826, 6.065066, 
    6.087969, 6.09293, 6.089534, 6.102671, 6.064328, 6.079013, 5.966931, 
    5.967578, 5.970622, 5.957223, 5.956419, 5.944223, 5.955099, 5.95971, 
    5.971514, 5.978412, 5.984989, 5.999462, 6.015565, 6.03818, 6.056235, 
    6.067171, 6.060482, 6.066385, 6.059776, 6.05669, 6.091054, 6.071726, 
    6.10078, 6.099181, 6.086006, 6.099362, 5.968038, 5.964302, 5.951252, 
    5.961465, 5.942899, 5.953256, 5.959194, 5.982192, 5.987295, 5.991948, 
    6.001197, 6.013024, 6.033774, 6.053636, 6.07024, 6.069028, 6.069453, 
    6.073138, 6.063975, 6.074646, 6.076412, 6.071754, 6.098965, 6.09119, 
    6.099146, 6.09409, 5.965523, 5.971808, 5.968414, 5.974776, 5.970279, 
    5.99021, 5.996189, 6.02422, 6.012777, 6.031063, 6.014654, 6.017546, 
    6.03155, 6.015557, 6.052585, 6.026816, 6.073282, 6.047391, 6.07479, 
    6.070168, 6.077847, 6.084699, 6.09337, 6.109308, 6.105626, 6.119005, 
    5.981166, 5.989267, 5.988602, 5.997118, 6.0034, 6.017075, 6.038968, 
    6.030749, 6.045895, 6.04892, 6.025939, 6.039999, 5.994728, 6.001993, 
    5.997705, 5.981777, 6.032577, 6.006477, 6.056496, 6.040595, 6.083715, 
    6.06307, 6.103589, 6.120813, 6.137269, 6.156254, 5.993743, 5.988231, 
    5.998145, 6.011757, 6.024531, 6.041448, 6.043206, 6.046363, 6.056356, 
    6.06327, 6.047315, 6.065009, 6.00358, 6.034865, 5.986103, 6.000726, 
    6.010976, 6.006529, 6.029822, 6.035297, 6.059307, 6.046072, 6.116518, 
    6.086078, 6.170887, 6.14711, 5.986294, 5.993747, 6.0196, 6.007308, 
    6.042603, 6.053029, 6.060135, 6.069144, 6.070152, 6.0755, 6.066732, 
    6.075173, 6.041484, 6.0575, 6.016702, 6.02617, 6.021831, 6.017035, 
    6.031831, 6.047526, 6.04794, 6.054713, 6.068748, 6.042748, 6.120306, 
    6.073303, 6.001867, 6.016104, 6.018233, 6.012699, 6.050408, 6.036726, 
    6.075381, 6.06541, 6.081771, 6.073632, 6.072431, 6.062003, 6.055494, 
    6.037338, 6.024025, 6.013511, 6.015961, 6.027514, 6.048505, 6.070209, 
    6.065824, 6.080528, 6.040039, 6.057973, 6.049939, 6.068099, 6.030513, 
    6.062535, 6.022757, 6.026104, 6.036456, 6.059021, 6.063748, 6.068658, 
    6.065644, 6.049053, 6.046659, 6.036223, 6.033305, 6.025381, 6.018786, 
    6.024792, 6.031085, 6.049091, 6.067054, 6.084785, 6.089157, 6.109705, 
    6.092868, 6.120552, 6.096849, 6.137984, 6.064407, 6.096312, 6.036953, 
    6.043163, 6.056071, 6.081882, 6.068023, 6.08427, 6.046571, 6.027874, 
    6.023135, 6.014136, 6.02334, 6.022595, 6.031401, 6.028575, 6.049691, 
    6.038348, 6.07238, 6.084161, 6.117574, 6.138042, 6.159029, 6.168261, 
    6.171079, 6.172253 ;

 EFLX_LH_TOT_R =
  5.945704, 5.96459, 5.960935, 5.976095, 5.967731, 5.977613, 5.949567, 
    5.965309, 5.955278, 5.947451, 6.005329, 5.976777, 6.035303, 6.017036, 
    6.064812, 6.032414, 6.071017, 6.064003, 6.08531, 6.079208, 6.106329, 
    6.088128, 6.12053, 6.102022, 6.104887, 6.087515, 5.982594, 6.001753, 
    5.981442, 5.984177, 5.982967, 5.967877, 5.960184, 5.944315, 5.947209, 
    5.958894, 5.985409, 5.976478, 5.999142, 5.998631, 6.023797, 6.012445, 
    6.056595, 6.0428, 6.079464, 6.070662, 6.079037, 6.076507, 6.079071, 
    6.066167, 6.07169, 6.060366, 6.014556, 6.027471, 5.988921, 5.965604, 
    5.950243, 5.939291, 5.940838, 5.943774, 5.958961, 5.973293, 5.984146, 
    5.991398, 5.998557, 6.020007, 6.031534, 6.058997, 6.054414, 6.062228, 
    6.069789, 6.082406, 6.080338, 6.085884, 6.062068, 6.077869, 6.050041, 
    6.058909, 6.000245, 5.978899, 5.969609, 5.961628, 5.942023, 5.955546, 
    5.950208, 5.962965, 5.971028, 5.967055, 5.991597, 5.982049, 6.032218, 
    6.010608, 6.068908, 6.05536, 6.072166, 6.0636, 6.07826, 6.065066, 
    6.087969, 6.09293, 6.089534, 6.102671, 6.064328, 6.079013, 5.966931, 
    5.967578, 5.970622, 5.957223, 5.956419, 5.944223, 5.955099, 5.95971, 
    5.971514, 5.978412, 5.984989, 5.999462, 6.015565, 6.03818, 6.056235, 
    6.067171, 6.060482, 6.066385, 6.059776, 6.05669, 6.091054, 6.071726, 
    6.10078, 6.099181, 6.086006, 6.099362, 5.968038, 5.964302, 5.951252, 
    5.961465, 5.942899, 5.953256, 5.959194, 5.982192, 5.987295, 5.991948, 
    6.001197, 6.013024, 6.033774, 6.053636, 6.07024, 6.069028, 6.069453, 
    6.073138, 6.063975, 6.074646, 6.076412, 6.071754, 6.098965, 6.09119, 
    6.099146, 6.09409, 5.965523, 5.971808, 5.968414, 5.974776, 5.970279, 
    5.99021, 5.996189, 6.02422, 6.012777, 6.031063, 6.014654, 6.017546, 
    6.03155, 6.015557, 6.052585, 6.026816, 6.073282, 6.047391, 6.07479, 
    6.070168, 6.077847, 6.084699, 6.09337, 6.109308, 6.105626, 6.119005, 
    5.981166, 5.989267, 5.988602, 5.997118, 6.0034, 6.017075, 6.038968, 
    6.030749, 6.045895, 6.04892, 6.025939, 6.039999, 5.994728, 6.001993, 
    5.997705, 5.981777, 6.032577, 6.006477, 6.056496, 6.040595, 6.083715, 
    6.06307, 6.103589, 6.120813, 6.137269, 6.156254, 5.993743, 5.988231, 
    5.998145, 6.011757, 6.024531, 6.041448, 6.043206, 6.046363, 6.056356, 
    6.06327, 6.047315, 6.065009, 6.00358, 6.034865, 5.986103, 6.000726, 
    6.010976, 6.006529, 6.029822, 6.035297, 6.059307, 6.046072, 6.116518, 
    6.086078, 6.170887, 6.14711, 5.986294, 5.993747, 6.0196, 6.007308, 
    6.042603, 6.053029, 6.060135, 6.069144, 6.070152, 6.0755, 6.066732, 
    6.075173, 6.041484, 6.0575, 6.016702, 6.02617, 6.021831, 6.017035, 
    6.031831, 6.047526, 6.04794, 6.054713, 6.068748, 6.042748, 6.120306, 
    6.073303, 6.001867, 6.016104, 6.018233, 6.012699, 6.050408, 6.036726, 
    6.075381, 6.06541, 6.081771, 6.073632, 6.072431, 6.062003, 6.055494, 
    6.037338, 6.024025, 6.013511, 6.015961, 6.027514, 6.048505, 6.070209, 
    6.065824, 6.080528, 6.040039, 6.057973, 6.049939, 6.068099, 6.030513, 
    6.062535, 6.022757, 6.026104, 6.036456, 6.059021, 6.063748, 6.068658, 
    6.065644, 6.049053, 6.046659, 6.036223, 6.033305, 6.025381, 6.018786, 
    6.024792, 6.031085, 6.049091, 6.067054, 6.084785, 6.089157, 6.109705, 
    6.092868, 6.120552, 6.096849, 6.137984, 6.064407, 6.096312, 6.036953, 
    6.043163, 6.056071, 6.081882, 6.068023, 6.08427, 6.046571, 6.027874, 
    6.023135, 6.014136, 6.02334, 6.022595, 6.031401, 6.028575, 6.049691, 
    6.038348, 6.07238, 6.084161, 6.117574, 6.138042, 6.159029, 6.168261, 
    6.171079, 6.172253 ;

 EFLX_LH_TOT_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 ELAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 ER =
  6.35757e-08, 6.385525e-08, 6.38009e-08, 6.402639e-08, 6.39013e-08, 
    6.404895e-08, 6.363237e-08, 6.386636e-08, 6.371699e-08, 6.360087e-08, 
    6.446398e-08, 6.403645e-08, 6.490803e-08, 6.463537e-08, 6.532027e-08, 
    6.48656e-08, 6.541195e-08, 6.530715e-08, 6.562256e-08, 6.55322e-08, 
    6.593564e-08, 6.566426e-08, 6.614476e-08, 6.587083e-08, 6.591368e-08, 
    6.565531e-08, 6.412248e-08, 6.441076e-08, 6.41054e-08, 6.41465e-08, 
    6.412806e-08, 6.390389e-08, 6.379094e-08, 6.355432e-08, 6.359728e-08, 
    6.377105e-08, 6.416499e-08, 6.403126e-08, 6.436827e-08, 6.436066e-08, 
    6.473585e-08, 6.456669e-08, 6.519728e-08, 6.501806e-08, 6.553597e-08, 
    6.540572e-08, 6.552985e-08, 6.549221e-08, 6.553034e-08, 6.533932e-08, 
    6.542116e-08, 6.525307e-08, 6.459837e-08, 6.479079e-08, 6.421691e-08, 
    6.387185e-08, 6.364264e-08, 6.347999e-08, 6.350298e-08, 6.354682e-08, 
    6.377208e-08, 6.398385e-08, 6.414524e-08, 6.42532e-08, 6.435957e-08, 
    6.468156e-08, 6.485197e-08, 6.523354e-08, 6.516466e-08, 6.528133e-08, 
    6.539276e-08, 6.557987e-08, 6.554907e-08, 6.563151e-08, 6.527824e-08, 
    6.551303e-08, 6.512544e-08, 6.523145e-08, 6.438852e-08, 6.406734e-08, 
    6.393085e-08, 6.381136e-08, 6.352067e-08, 6.372141e-08, 6.364228e-08, 
    6.383054e-08, 6.395017e-08, 6.3891e-08, 6.425615e-08, 6.411419e-08, 
    6.486207e-08, 6.453993e-08, 6.537977e-08, 6.51788e-08, 6.542793e-08, 
    6.53008e-08, 6.551863e-08, 6.532259e-08, 6.566219e-08, 6.573613e-08, 
    6.56856e-08, 6.587971e-08, 6.531172e-08, 6.552985e-08, 6.388935e-08, 
    6.389899e-08, 6.394394e-08, 6.374634e-08, 6.373425e-08, 6.355315e-08, 
    6.371429e-08, 6.378291e-08, 6.39571e-08, 6.406013e-08, 6.415808e-08, 
    6.437342e-08, 6.461393e-08, 6.495023e-08, 6.519183e-08, 6.535377e-08, 
    6.525447e-08, 6.534214e-08, 6.524414e-08, 6.519819e-08, 6.570843e-08, 
    6.542193e-08, 6.585179e-08, 6.5828e-08, 6.563347e-08, 6.583068e-08, 
    6.390577e-08, 6.385024e-08, 6.365745e-08, 6.380832e-08, 6.353343e-08, 
    6.36873e-08, 6.377579e-08, 6.411717e-08, 6.419216e-08, 6.426171e-08, 
    6.439907e-08, 6.457535e-08, 6.488458e-08, 6.515364e-08, 6.539925e-08, 
    6.538125e-08, 6.538759e-08, 6.544246e-08, 6.530654e-08, 6.546477e-08, 
    6.549133e-08, 6.542189e-08, 6.582482e-08, 6.570971e-08, 6.58275e-08, 
    6.575254e-08, 6.386828e-08, 6.396172e-08, 6.391124e-08, 6.400618e-08, 
    6.393929e-08, 6.423671e-08, 6.432588e-08, 6.474312e-08, 6.457188e-08, 
    6.484441e-08, 6.459956e-08, 6.464295e-08, 6.485331e-08, 6.461279e-08, 
    6.513881e-08, 6.47822e-08, 6.544459e-08, 6.508849e-08, 6.546691e-08, 
    6.539818e-08, 6.551196e-08, 6.561386e-08, 6.574206e-08, 6.59786e-08, 
    6.592382e-08, 6.612164e-08, 6.410102e-08, 6.422221e-08, 6.421153e-08, 
    6.433836e-08, 6.443215e-08, 6.463544e-08, 6.496149e-08, 6.483888e-08, 
    6.506396e-08, 6.510916e-08, 6.476719e-08, 6.497716e-08, 6.430331e-08, 
    6.441219e-08, 6.434736e-08, 6.411058e-08, 6.486714e-08, 6.447888e-08, 
    6.519582e-08, 6.498549e-08, 6.559934e-08, 6.529407e-08, 6.589367e-08, 
    6.615002e-08, 6.639124e-08, 6.667317e-08, 6.428834e-08, 6.4206e-08, 
    6.435344e-08, 6.455743e-08, 6.47467e-08, 6.499832e-08, 6.502406e-08, 
    6.507121e-08, 6.51933e-08, 6.529596e-08, 6.508611e-08, 6.53217e-08, 
    6.443745e-08, 6.490084e-08, 6.417487e-08, 6.439348e-08, 6.454541e-08, 
    6.447876e-08, 6.482487e-08, 6.490644e-08, 6.523793e-08, 6.506657e-08, 
    6.608675e-08, 6.56354e-08, 6.688783e-08, 6.653783e-08, 6.417723e-08, 
    6.428806e-08, 6.467379e-08, 6.449026e-08, 6.501512e-08, 6.514431e-08, 
    6.524932e-08, 6.538358e-08, 6.539807e-08, 6.547761e-08, 6.534727e-08, 
    6.547247e-08, 6.499886e-08, 6.52105e-08, 6.46297e-08, 6.477106e-08, 
    6.470603e-08, 6.463469e-08, 6.485485e-08, 6.508942e-08, 6.509442e-08, 
    6.516963e-08, 6.53816e-08, 6.501724e-08, 6.614502e-08, 6.544855e-08, 
    6.440892e-08, 6.462241e-08, 6.465289e-08, 6.457019e-08, 6.513136e-08, 
    6.492802e-08, 6.547567e-08, 6.532767e-08, 6.557018e-08, 6.544967e-08, 
    6.543194e-08, 6.527716e-08, 6.51808e-08, 6.493735e-08, 6.473926e-08, 
    6.458218e-08, 6.46187e-08, 6.479126e-08, 6.510376e-08, 6.539939e-08, 
    6.533463e-08, 6.555175e-08, 6.497706e-08, 6.521804e-08, 6.512491e-08, 
    6.536776e-08, 6.483562e-08, 6.528879e-08, 6.471979e-08, 6.476968e-08, 
    6.492399e-08, 6.52344e-08, 6.530306e-08, 6.537638e-08, 6.533113e-08, 
    6.51117e-08, 6.507574e-08, 6.492024e-08, 6.487731e-08, 6.475882e-08, 
    6.466072e-08, 6.475035e-08, 6.484448e-08, 6.511178e-08, 6.535268e-08, 
    6.561532e-08, 6.567959e-08, 6.598647e-08, 6.573666e-08, 6.61489e-08, 
    6.579844e-08, 6.64051e-08, 6.531504e-08, 6.578811e-08, 6.493101e-08, 
    6.502334e-08, 6.519036e-08, 6.557342e-08, 6.536661e-08, 6.560847e-08, 
    6.507433e-08, 6.479721e-08, 6.47255e-08, 6.459173e-08, 6.472857e-08, 
    6.471743e-08, 6.484837e-08, 6.480629e-08, 6.512066e-08, 6.49518e-08, 
    6.54315e-08, 6.560656e-08, 6.610091e-08, 6.640397e-08, 6.671245e-08, 
    6.684864e-08, 6.689009e-08, 6.690742e-08 ;

 ERRH2O =
  -22839, -22872.79, -22866.16, -22893.82, -22878.42, -22896.62, -22845.79, 
    -22874.14, -22855.99, -22842.01, -22948.74, -22895.07, -23006.17, 
    -22970.66, -23060.56, -23000.59, -23072.89, -23058.81, -23101.57, 
    -23089.2, -23145.18, -23107.31, -23175.03, -23136.05, -23142.08, 
    -23106.07, -22905.75, -22941.99, -22903.63, -22908.75, -22906.45, 
    -22878.74, -22864.95, -22836.44, -22841.58, -22862.54, -22911.06, 
    -22894.42, -22936.61, -22935.65, -22983.65, -22961.84, -23044.18, 
    -23020.62, -23089.72, -23072.05, -23088.88, -23083.76, -23088.95, 
    -23063.12, -23074.13, -23051.59, -22965.9, -22990.8, -22917.57, 
    -22874.82, -22847.02, -22827.58, -22830.32, -22835.54, -22862.66, 
    -22888.57, -22908.59, -22922.13, -22935.51, -22976.62, -22998.8, 
    -23048.99, -23039.87, -23055.36, -23070.3, -23095.72, -23091.51, 
    -23102.8, -23054.94, -23086.59, -23034.69, -23048.71, -22939.18, 
    -22898.9, -22882.05, -22867.43, -22832.42, -22856.52, -22846.98, 
    -22869.77, -22884.42, -22877.16, -22922.5, -22904.72, -23000.13, 
    -22958.41, -23068.55, -23041.73, -23075.04, -23057.96, -23087.36, 
    -23060.87, -23107.02, -23117.25, -23110.25, -23137.3, -23059.42, 
    -23088.88, -22876.95, -22878.14, -22883.65, -22859.54, -22858.07, 
    -22836.3, -22855.66, -22863.97, -22885.27, -22898, -22910.2, -22937.26, 
    -22967.9, -23011.73, -23043.46, -23065.05, -23051.78, -23063.49, 
    -23050.4, -23044.3, -23113.41, -23074.23, -23133.38, -23130.04, 
    -23103.07, -23130.42, -22878.97, -22872.17, -22848.8, -22867.06, 
    -22833.95, -22852.4, -22863.11, -22905.09, -22914.46, -22923.2, -22940.5, 
    -22962.95, -23003.08, -23038.41, -23071.17, -23068.75, -23069.6, 
    -23077.01, -23058.72, -23080.03, -23083.64, -23074.23, -23129.6, 
    -23113.58, -23129.97, -23119.53, -22874.38, -22885.84, -22879.64, 
    -22891.32, -22883.08, -22920.05, -22931.27, -22984.6, -22962.5, 
    -22997.81, -22966.05, -22971.64, -22998.98, -22967.75, -23036.46, 
    -22989.68, -23077.3, -23029.84, -23080.32, -23071.03, -23086.45, 
    -23100.38, -23118.07, -23151.26, -23143.51, -23171.7, -22903.08, 
    -22918.23, -22916.89, -22932.84, -22944.69, -22970.67, -23013.22, 
    -22997.09, -23026.62, -23032.55, -22987.73, -23015.29, -22928.43, 
    -22942.17, -22933.97, -22904.27, -23000.79, -22950.63, -23043.99, 
    -23016.37, -23098.38, -23057.06, -23139.26, -23175.79, -23210.88, 
    -23252.65, -22926.55, -22916.2, -22934.74, -22960.65, -22985.06, 
    -23018.04, -23021.4, -23027.56, -23043.65, -23057.31, -23029.52, 
    -23060.75, -22945.37, -23005.22, -22912.3, -22939.8, -22959.11, 
    -22950.61, -22995.25, -23005.96, -23049.58, -23026.96, -23166.69, 
    -23103.34, -23284.78, -23232.62, -22912.59, -22926.52, -22975.62, 
    -22952.07, -23020.23, -23037.18, -23051.09, -23069.06, -23071.01, 
    -23081.78, -23064.18, -23081.08, -23018.11, -23045.93, -22969.93, 
    -22988.23, -22979.79, -22970.57, -22999.18, -23029.96, -23030.61, 
    -23040.52, -23068.8, -23020.51, -23175.07, -23077.84, -22941.75, 
    -22968.99, -22972.92, -22962.28, -23035.47, -23008.8, -23081.51, 
    -23061.55, -23094.39, -23077.99, -23075.59, -23054.8, -23042, -23010.03, 
    -22984.1, -22963.82, -22968.51, -22990.86, -23031.84, -23071.19, 
    -23062.49, -23091.87, -23015.27, -23046.93, -23034.62, -23066.93, 
    -22996.66, -23056.36, -22981.57, -22988.05, -23008.27, -23049.11, 
    -23058.26, -23068.09, -23062.02, -23032.88, -23028.16, -23007.77, 
    -23002.12, -22986.64, -22973.93, -22985.54, -22997.82, -23032.89, 
    -23064.91, -23100.58, -23109.42, -23152.38, -23117.32, -23175.63, 
    -23125.93, -23212.92, -23059.87, -23124.48, -23009.2, -23021.3, 
    -23043.27, -23094.84, -23066.78, -23099.64, -23027.97, -22991.64, 
    -22982.31, -22965.05, -22982.71, -22981.26, -22998.33, -22992.82, 
    -23034.06, -23011.94, -23075.53, -23099.38, -23168.72, -23212.75, 
    -23258.49, -23278.87, -23285.12, -23287.74 ;

 ERRH2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ERRSEB =
  -5.554146e-15, -8.368608e-15, -1.097268e-14, -1.020937e-14, -1.035655e-15, 
    -9.835425e-15, -2.989683e-15, -1.267431e-14, -4.876899e-15, 
    -8.687409e-15, -7.671896e-15, -9.205839e-15, -1.072132e-14, 
    -6.272696e-16, 2.44316e-15, 2.546362e-16, -1.625905e-14, -5.469636e-15, 
    2.796913e-15, -1.42854e-14, -2.290752e-15, -1.47739e-14, -5.16156e-15, 
    -3.092677e-15, -1.611659e-14, -1.457792e-14, -7.643099e-15, 
    -6.660791e-15, -1.0229e-14, -4.828733e-16, -9.401195e-15, -2.124881e-15, 
    -1.46414e-14, -9.908645e-15, -3.337258e-15, -3.210523e-15, -1.703362e-14, 
    -1.362275e-14, -1.139102e-14, -1.32119e-14, -1.022889e-14, -9.14119e-15, 
    -1.182459e-14, -1.159211e-14, -1.383656e-14, -1.005241e-14, 1.505029e-15, 
    -1.063174e-14, -8.685157e-15, -1.575019e-14, -1.445188e-14, 
    -4.224352e-15, -7.916475e-15, -6.662718e-15, -8.966172e-15, -9.81658e-15, 
    5.871755e-15, 5.144418e-16, -1.493527e-14, -8.974621e-15, -1.887772e-15, 
    -2.662461e-15, -1.018665e-14, -8.396308e-15, -5.515037e-15, 
    -4.631344e-15, -1.133774e-14, 4.110537e-15, -1.302756e-14, -1.171064e-14, 
    -1.507879e-14, -9.308696e-15, -1.172846e-14, -9.461339e-15, 
    -1.360633e-14, -1.862076e-14, -1.529667e-14, -9.73903e-15, -8.85861e-15, 
    -1.136495e-14, -5.465744e-15, 1.208162e-15, -1.136831e-14, -1.834613e-14, 
    -5.96674e-15, -1.314833e-14, -9.736146e-15, -3.112514e-15, -6.98441e-15, 
    -1.307466e-14, -1.603653e-15, -1.316161e-14, -1.010746e-14, 
    -1.258644e-14, -1.603832e-14, -1.120563e-14, -6.374222e-15, 3.323624e-16, 
    -1.13889e-14, -8.137849e-15, -1.324221e-14, -1.266395e-14, -1.23415e-14, 
    -5.07393e-15, -6.364192e-15, -1.387557e-14, -9.361944e-15, -5.638916e-15, 
    -1.074755e-14, -1.066911e-14, -1.060444e-14, -1.158943e-14, -7.8955e-16, 
    -1.041486e-14, -8.029981e-15, -1.445913e-15, -6.973067e-15, 
    -6.324666e-15, -8.858913e-15, -1.163813e-14, -5.565525e-15, -3.25699e-15, 
    -1.292843e-14, -1.131602e-14, -8.509208e-15, 1.928536e-16, 2.057208e-15, 
    -7.446517e-15, -1.566144e-15, -1.41475e-14, -1.157924e-14, -6.464217e-15, 
    -9.97369e-15, -6.3062e-15, -5.110233e-15, -2.452283e-14, -1.159035e-14, 
    -1.01002e-14, -2.934837e-15, -3.67197e-15, -1.74723e-14, -7.791069e-15, 
    -1.356388e-14, -1.054131e-14, -6.403537e-15, -7.964066e-15, 
    -1.276227e-14, -3.622419e-15, -2.565554e-15, -7.871847e-15, 
    -1.075355e-14, -1.071449e-14, -9.072144e-15, -1.414558e-14, 
    -1.145442e-14, -4.939216e-15, -1.319198e-14, -2.019073e-15, 
    -2.325371e-15, -2.33502e-15, -3.060052e-15, -8.722537e-15, -5.307292e-15, 
    -1.290579e-14, -3.174736e-15, -1.047885e-14, -8.748734e-15, 
    -1.235722e-14, 4.260978e-16, -2.004331e-14, -1.493468e-14, -9.164752e-15, 
    -7.791393e-15, -1.002516e-15, -1.695062e-14, -1.259635e-14, 
    -1.147301e-14, -1.235158e-15, 1.770354e-16, -9.341709e-15, -6.985997e-15, 
    1.256477e-15, 9.677259e-17, -3.998307e-15, -1.088368e-14, -3.27363e-15, 
    -1.424211e-14, -3.681609e-15, -1.58474e-14, -7.03253e-15, -4.137834e-15, 
    -9.988024e-15, -7.319427e-15, -4.238363e-15, -1.22346e-14, -6.201269e-15, 
    -1.121877e-14, -8.471602e-16, -1.388261e-14, -9.127057e-15, 
    -1.556236e-15, -4.386866e-15, -8.323809e-15, -9.02591e-15, -6.427307e-15, 
    -3.96786e-15, -1.367968e-14, -2.165459e-15, -1.186672e-14, -1.323497e-14, 
    8.847888e-16, -3.480716e-15, -6.441088e-15, -1.569754e-14, -6.172863e-15, 
    -1.677447e-14, -1.417032e-15, -6.817553e-15, -6.971583e-15, -1.20509e-14, 
    -9.094389e-15, -1.481575e-14, -3.639063e-16, -1.890243e-14, 
    -7.077695e-15, -1.899361e-14, -1.046081e-14, -1.265931e-15, 
    -1.429673e-14, -7.630985e-15, -1.691088e-14, -1.194523e-14, 
    -9.148882e-15, -1.063519e-14, -1.402115e-14, -6.552476e-15, 
    -6.060709e-15, -2.045772e-15, -3.243504e-15, -9.677406e-15, -5.5231e-15, 
    -7.971412e-15, -7.7241e-16, -2.104353e-15, -2.465534e-14, -9.708482e-15, 
    -1.277822e-14, -7.969702e-15, -1.23402e-15, -8.232026e-15, -5.124367e-15, 
    -1.797933e-14, -6.461989e-15, -1.958821e-15, -9.596874e-15, 
    -1.323989e-14, -7.578954e-15, -9.375573e-15, -7.258524e-15, 
    -2.650185e-15, -1.39916e-14, -1.09776e-14, -8.598757e-15, -8.539951e-15, 
    -3.378321e-15, -4.682942e-15, -1.735452e-14, -1.309574e-14, 
    -8.427873e-15, -7.067095e-15, -8.695578e-15, -1.260191e-14, 
    -8.216535e-15, -1.346902e-14, -1.204486e-14, -7.864592e-15, 
    -7.916865e-15, -2.225829e-14, -1.286198e-14, -1.371396e-15, -2.32532e-15, 
    -2.581973e-15, -1.594607e-14, -1.833325e-14, -1.401912e-14, 
    -1.885682e-14, -9.411565e-15, -7.727202e-15, -8.998883e-15, 
    -1.515049e-14, -1.697176e-14, -7.574707e-15, -7.705452e-15, -4.21654e-15, 
    -1.029189e-14, -5.198778e-15, -1.410067e-14, -1.924429e-15, 
    -5.237513e-16, -8.342046e-15, -5.00272e-15, -8.060172e-15, -9.828077e-15, 
    -8.130987e-15, -8.666175e-15, -9.194405e-15, -1.433115e-14, 
    -1.220201e-14, -1.18861e-14, -1.102274e-14, -6.527695e-15, -5.178767e-15, 
    -1.666952e-14, -9.82373e-15, -1.693432e-14, -1.501693e-14, -8.616626e-15, 
    8.557158e-16, -6.773058e-15, -1.273825e-14, -1.339711e-14, -5.901013e-15, 
    -9.66003e-15, -1.52956e-14, -3.849817e-15, -3.1595e-15, -1.121501e-14, 
    -1.666213e-15, -1.310606e-14, -1.095282e-14, -1.145955e-14, 
    -1.037719e-14, -7.871213e-15, -1.814287e-14, -5.315795e-15, 
    -7.946584e-15, -1.122492e-14, -1.247093e-14 ;

 ERRSOI =
  -3.055317e-10, -2.413545e-10, -2.661513e-10, -3.10494e-10, -2.15602e-10, 
    -3.295109e-10, -3.064284e-10, -2.312958e-10, -3.501749e-10, 
    -3.228471e-10, -3.435995e-10, -2.582257e-10, -3.061282e-10, 
    -2.000983e-10, -4.173785e-10, -2.727582e-10, -2.618215e-10, 
    -3.256279e-10, -3.781273e-10, -2.827255e-10, -2.126646e-10, 
    -3.192806e-11, -2.365083e-10, -4.79105e-10, -3.26496e-10, -1.822068e-10, 
    -1.439647e-10, -2.719009e-10, -1.930931e-10, -3.810874e-10, 
    -2.314239e-10, -2.458453e-10, -3.728499e-10, -4.199934e-10, 
    -3.411334e-10, -3.209266e-10, -3.168557e-10, -4.366163e-10, 
    -4.719954e-10, -2.429944e-10, 4.813402e-11, -3.594098e-10, -2.293907e-10, 
    -4.850168e-10, -2.739475e-10, -2.974825e-10, -3.243553e-10, 
    -1.827325e-10, -1.065222e-10, -1.560447e-10, -3.106775e-10, -3.84672e-10, 
    -2.809735e-10, -8.326662e-11, -4.027662e-10, -2.550594e-10, 
    -3.392643e-10, -2.901509e-10, -3.722864e-10, -3.8265e-10, -2.808625e-10, 
    -2.067775e-10, -3.378181e-10, -3.154309e-10, -3.22483e-10, -2.177839e-10, 
    -4.060912e-10, -1.287238e-10, -3.65773e-10, -5.057217e-10, -1.488821e-10, 
    -3.810319e-10, -3.660245e-10, -4.22786e-10, -4.690039e-10, -3.604563e-10, 
    -2.356644e-10, -2.607869e-10, -2.278809e-10, -3.436798e-10, 
    -3.946687e-10, -1.909077e-10, -5.332635e-10, -3.226663e-10, 
    -2.516798e-10, -2.686939e-10, -1.737693e-10, -4.178439e-10, 
    -2.592496e-10, -2.481534e-10, -2.322194e-10, -4.365465e-10, 
    -3.432706e-10, -2.782435e-10, -2.452418e-10, -4.045231e-10, 
    -2.152074e-10, -3.021282e-10, -2.295767e-10, -2.418445e-10, 
    -1.970306e-10, -3.433437e-10, -3.168475e-10, -2.821508e-10, 
    -3.376794e-10, -3.963874e-10, -2.271662e-10, -2.522767e-10, 
    -4.278939e-10, -2.39706e-10, -2.321656e-10, -2.584863e-10, -4.271115e-10, 
    -4.090446e-10, -2.770204e-10, -3.46296e-10, -2.806335e-10, -3.026688e-10, 
    -4.932959e-10, -3.667982e-10, -2.236086e-10, -1.958223e-10, 
    -1.997918e-10, -4.213171e-10, -2.98049e-10, -1.062737e-10, -2.757374e-10, 
    -1.109269e-10, -1.273952e-10, -2.093272e-10, -3.683182e-10, 
    -3.064884e-11, -1.661085e-10, -3.620242e-10, -4.023815e-10, 
    -3.101457e-10, -1.981268e-10, -2.280585e-10, -1.195248e-10, 
    -4.021628e-10, -3.211966e-10, -3.852614e-10, -2.878211e-10, 
    -3.674166e-10, -2.108393e-10, -2.256748e-10, -3.422787e-10, -2.75291e-10, 
    -3.122602e-10, -2.407452e-10, -2.497408e-10, -2.751446e-10, 
    -2.915387e-10, -2.814835e-10, -9.127369e-11, -3.860731e-10, 
    -2.400132e-10, -3.48557e-10, -4.107113e-10, -2.918315e-10, -1.063249e-10, 
    -3.553663e-10, -5.053414e-10, -2.829545e-10, -2.417782e-10, 
    -4.775503e-10, -3.16045e-10, -1.41416e-10, -4.069514e-10, -1.156109e-10, 
    -2.734528e-10, -2.041609e-10, -3.151392e-10, -2.918768e-10, 
    -1.579964e-10, -1.989471e-10, -3.706551e-10, -3.010041e-10, 
    -4.890552e-10, -1.871386e-10, -3.363674e-10, -4.406318e-10, -1.7287e-10, 
    -3.112437e-10, -3.925991e-10, -2.919568e-10, -4.553808e-10, 
    -4.392058e-10, -3.207399e-10, -1.29755e-10, -3.229953e-10, -5.381481e-10, 
    -2.692205e-10, -2.947161e-10, -3.156067e-10, -3.418533e-10, 
    -1.419738e-10, -2.275911e-10, -3.212705e-10, -3.710059e-10, 
    -1.350115e-10, -2.08513e-10, -2.441814e-10, -2.918128e-10, -2.95174e-10, 
    -2.654728e-10, -1.565299e-10, -1.986181e-10, -2.754137e-10, 
    -3.962219e-10, -2.596777e-10, -1.780508e-10, -1.251112e-10, 
    -4.724856e-11, -2.554988e-10, -2.686445e-10, -3.001691e-10, 
    -4.157256e-10, -3.919963e-10, -1.843041e-10, -2.254959e-10, 
    -3.106976e-10, -2.448081e-10, -3.942349e-10, -3.413587e-10, 
    -1.826665e-10, -2.101508e-10, -3.220086e-10, -3.097902e-10, 
    -2.404569e-10, -1.746224e-10, -3.543465e-10, -1.664652e-10, 
    -3.616436e-10, -2.523853e-10, -5.488524e-10, -2.649112e-10, 
    -2.734261e-10, -2.413089e-10, -4.280974e-10, -4.972271e-10, 
    -3.791374e-10, -2.590499e-10, -4.955611e-10, -2.395755e-10, 
    -3.702062e-10, -3.836838e-10, -2.427963e-10, -1.743265e-10, 
    -3.921988e-10, -8.072861e-11, -3.440209e-10, -3.289062e-10, 
    -3.804906e-10, -4.261101e-10, -2.647388e-10, -3.517685e-10, 
    -1.840527e-10, -1.885059e-10, -1.245408e-10, -4.144959e-10, 
    -2.393683e-10, -4.59147e-10, -2.703301e-10, -1.835832e-10, -2.271528e-10, 
    -2.305254e-10, -3.687458e-10, -3.497909e-10, -3.621681e-10, 
    -2.903134e-10, -5.071654e-10, -1.825396e-10, -3.688373e-10, 
    -1.775101e-10, -2.49079e-10, -3.715161e-10, -4.055452e-10, -5.321824e-10, 
    -2.331774e-10, -3.461281e-10, -2.417869e-10, -3.863279e-10, 
    -2.452077e-10, -5.216905e-10, -3.381993e-10, -2.044867e-10, 
    -5.090913e-10, -2.597786e-10, -6.042506e-11, -1.261945e-10, 
    -3.321359e-10, -4.286475e-10, -1.984971e-10, -4.392e-10, -3.407405e-10, 
    -1.604557e-10, -3.028688e-10, -1.45157e-10, -3.081216e-10, -5.681949e-10, 
    -2.371157e-10, -1.178525e-10, -4.856066e-10, -1.054971e-10, 
    -3.566923e-10, -2.655402e-10, -3.176114e-10, -2.350545e-10, 
    -3.059828e-10, -2.102245e-10, -2.310328e-10, -2.180421e-10, 
    -3.243611e-10, -3.669587e-10, -2.803714e-10, -3.655026e-10, 
    -2.974667e-10, -3.032251e-10, -3.586493e-10, -2.825933e-10, 
    -2.041947e-10, -1.985599e-10, -2.093165e-10, -3.049831e-10, 
    -2.512947e-10, -3.128598e-10, -1.935881e-10, -2.694948e-10, 
    -3.228811e-10, -1.742828e-10, -4.560634e-10, -3.575615e-10, -3.14816e-10, 
    -1.649339e-10, -2.209107e-10, -3.85744e-10, -3.167429e-10 ;

 ERRSOL =
  1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17 ;

 ESAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 FAREA_BURNED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCEV =
  -1.621223, -1.620124, -1.620332, -1.619455, -1.619934, -1.619365, -1.62099, 
    -1.620089, -1.620659, -1.62111, -1.617776, -1.619413, -1.615986, 
    -1.617043, -1.614353, -1.616164, -1.613981, -1.614383, -1.613114, 
    -1.613477, -1.611894, -1.612946, -1.61103, -1.612133, -1.611969, 
    -1.612984, -1.619062, -1.617986, -1.619131, -1.618977, -1.619041, 
    -1.619932, -1.620394, -1.621291, -1.621125, -1.620457, -1.618906, 
    -1.619419, -1.61808, -1.61811, -1.616644, -1.617306, -1.614821, 
    -1.615521, -1.613461, -1.613986, -1.61349, -1.613637, -1.613488, 
    -1.614256, -1.613928, -1.614595, -1.617187, -1.616433, -1.618694, 
    -1.620089, -1.620955, -1.621584, -1.621496, -1.621331, -1.620454, 
    -1.619606, -1.618965, -1.618539, -1.618115, -1.616901, -1.616207, 
    -1.614689, -1.614945, -1.614496, -1.614037, -1.613292, -1.613411, 
    -1.613087, -1.614493, -1.613567, -1.615091, -1.614681, -1.618078, 
    -1.619277, -1.619852, -1.620295, -1.621429, -1.620651, -1.62096, 
    -1.620208, -1.61974, -1.619968, -1.618527, -1.619092, -1.616166, 
    -1.617424, -1.61409, -1.614891, -1.613895, -1.6144, -1.613541, -1.614314, 
    -1.61296, -1.612672, -1.61287, -1.612082, -1.614359, -1.613497, 
    -1.619978, -1.619941, -1.619761, -1.620554, -1.620598, -1.6213, 
    -1.620669, -1.620406, -1.619707, -1.619307, -1.61892, -1.618068, 
    -1.617136, -1.615807, -1.61484, -1.614189, -1.614583, -1.614236, 
    -1.614627, -1.614807, -1.612785, -1.61393, -1.612196, -1.612289, 
    -1.613082, -1.612279, -1.619914, -1.620128, -1.620894, -1.620295, 
    -1.621375, -1.620781, -1.620444, -1.619097, -1.618781, -1.618512, 
    -1.617963, -1.617273, -1.616064, -1.615, -1.614007, -1.614078, -1.614054, 
    -1.61384, -1.614381, -1.61375, -1.613651, -1.613921, -1.612302, 
    -1.612765, -1.612292, -1.612591, -1.620057, -1.619693, -1.619891, 
    -1.619523, -1.619789, -1.618628, -1.618279, -1.616635, -1.617291, 
    -1.616225, -1.617177, -1.617013, -1.616224, -1.61712, -1.615074, 
    -1.61649, -1.613831, -1.615286, -1.613741, -1.614012, -1.613556, 
    -1.613156, -1.612637, -1.611698, -1.611912, -1.611112, -1.619143, 
    -1.618676, -1.618703, -1.618203, -1.617838, -1.617033, -1.615753, 
    -1.61623, -1.615337, -1.615163, -1.61651, -1.615698, -1.618352, 
    -1.617937, -1.618173, -1.619115, -1.61614, -1.617673, -1.614827, 
    -1.615654, -1.613215, -1.61445, -1.612034, -1.61103, -1.610011, 
    -1.608896, -1.618405, -1.618724, -1.618139, -1.617363, -1.6166, 
    -1.615606, -1.615497, -1.615314, -1.614828, -1.614421, -1.615271, 
    -1.614317, -1.617871, -1.616, -1.618858, -1.618014, -1.617402, -1.617655, 
    -1.616281, -1.615961, -1.614667, -1.615327, -1.611291, -1.613092, 
    -1.607992, -1.60944, -1.618839, -1.618399, -1.616897, -1.617608, 
    -1.615532, -1.61503, -1.614604, -1.614082, -1.614014, -1.613702, 
    -1.614215, -1.613717, -1.615604, -1.614764, -1.617051, -1.616504, 
    -1.616751, -1.617032, -1.616164, -1.615261, -1.615218, -1.614936, 
    -1.614168, -1.615523, -1.611102, -1.613889, -1.617921, -1.617112, 
    -1.616968, -1.617287, -1.615077, -1.615883, -1.613706, -1.614294, 
    -1.613325, -1.613809, -1.613881, -1.614495, -1.614883, -1.61585, 
    -1.616631, -1.617238, -1.617095, -1.616428, -1.6152, -1.614019, 
    -1.614283, -1.613398, -1.615684, -1.614744, -1.615113, -1.614138, 
    -1.616248, -1.614525, -1.616696, -1.616501, -1.615898, -1.614696, 
    -1.614392, -1.61411, -1.61428, -1.615164, -1.615299, -1.615907, 
    -1.616086, -1.616542, -1.616929, -1.616581, -1.61622, -1.615154, 
    -1.614207, -1.613154, -1.612886, -1.611706, -1.6127, -1.611091, 
    -1.612509, -1.610023, -1.614389, -1.612502, -1.615863, -1.615498, 
    -1.614866, -1.613344, -1.614142, -1.613197, -1.615303, -1.616417, 
    -1.616675, -1.617205, -1.616663, -1.616706, -1.616188, -1.616353, 
    -1.615118, -1.615782, -1.613889, -1.613199, -1.611204, -1.609986, 
    -1.6087, -1.608143, -1.607971, -1.6079 ;

 FCH4 =
  1.82798e-13, 1.82745e-13, 1.827561e-13, 1.827074e-13, 1.827353e-13, 
    1.827022e-13, 1.82788e-13, 1.827427e-13, 1.827724e-13, 1.827936e-13, 
    1.825911e-13, 1.827051e-13, 1.824381e-13, 1.825367e-13, 1.812103e-13, 
    1.824544e-13, 1.812158e-13, 1.812093e-13, 1.812148e-13, 1.812176e-13, 
    1.811763e-13, 1.812123e-13, 1.811248e-13, 1.81188e-13, 1.811805e-13, 
    1.812129e-13, 1.826845e-13, 1.826069e-13, 1.826887e-13, 1.826786e-13, 
    1.826831e-13, 1.827347e-13, 1.82758e-13, 1.828016e-13, 1.827943e-13, 
    1.82762e-13, 1.826739e-13, 1.827063e-13, 1.826193e-13, 1.826215e-13, 
    1.825021e-13, 1.825592e-13, 1.811976e-13, 1.811682e-13, 1.812175e-13, 
    1.812156e-13, 1.812176e-13, 1.812177e-13, 1.812176e-13, 1.812118e-13, 
    1.812162e-13, 1.812041e-13, 1.825489e-13, 1.824824e-13, 1.826606e-13, 
    1.827415e-13, 1.827862e-13, 1.82814e-13, 1.828102e-13, 1.828029e-13, 
    1.827618e-13, 1.827172e-13, 1.826789e-13, 1.826511e-13, 1.826218e-13, 
    1.82521e-13, 1.824596e-13, 1.81202e-13, 1.811932e-13, 1.81207e-13, 
    1.81215e-13, 1.812165e-13, 1.812173e-13, 1.812143e-13, 1.812067e-13, 
    1.812177e-13, 1.811873e-13, 1.812017e-13, 1.826134e-13, 1.826979e-13, 
    1.827289e-13, 1.82754e-13, 1.828073e-13, 1.827716e-13, 1.827862e-13, 
    1.827501e-13, 1.827247e-13, 1.827375e-13, 1.826503e-13, 1.826866e-13, 
    1.824558e-13, 1.825677e-13, 1.812143e-13, 1.811951e-13, 1.812164e-13, 
    1.812088e-13, 1.812177e-13, 1.812105e-13, 1.812124e-13, 1.81206e-13, 
    1.812107e-13, 1.811866e-13, 1.812097e-13, 1.812176e-13, 1.827378e-13, 
    1.827358e-13, 1.827261e-13, 1.827668e-13, 1.827691e-13, 1.828018e-13, 
    1.827729e-13, 1.827597e-13, 1.827232e-13, 1.826996e-13, 1.826757e-13, 
    1.826178e-13, 1.825438e-13, 1.824215e-13, 1.811969e-13, 1.812128e-13, 
    1.812043e-13, 1.81212e-13, 1.812032e-13, 1.811977e-13, 1.812087e-13, 
    1.812162e-13, 1.811911e-13, 1.811947e-13, 1.812142e-13, 1.811943e-13, 
    1.827343e-13, 1.82746e-13, 1.827835e-13, 1.827546e-13, 1.828052e-13, 
    1.82778e-13, 1.82761e-13, 1.826858e-13, 1.82667e-13, 1.826488e-13, 
    1.826104e-13, 1.825564e-13, 1.824472e-13, 1.811916e-13, 1.812153e-13, 
    1.812144e-13, 1.812147e-13, 1.812169e-13, 1.812092e-13, 1.812174e-13, 
    1.812177e-13, 1.812162e-13, 1.811952e-13, 1.812086e-13, 1.811948e-13, 
    1.812043e-13, 1.827423e-13, 1.827221e-13, 1.827332e-13, 1.827121e-13, 
    1.827271e-13, 1.826554e-13, 1.826312e-13, 1.824995e-13, 1.825575e-13, 
    1.824625e-13, 1.825485e-13, 1.825342e-13, 1.824591e-13, 1.825442e-13, 
    1.811893e-13, 1.824855e-13, 1.812169e-13, 1.811811e-13, 1.812174e-13, 
    1.812152e-13, 1.812177e-13, 1.812152e-13, 1.812054e-13, 1.811675e-13, 
    1.811787e-13, 1.811315e-13, 1.826898e-13, 1.826592e-13, 1.82662e-13, 
    1.826278e-13, 1.826007e-13, 1.825367e-13, 1.82417e-13, 1.824646e-13, 
    1.811769e-13, 1.811847e-13, 1.82491e-13, 1.824107e-13, 1.826375e-13, 
    1.826065e-13, 1.826252e-13, 1.826874e-13, 1.824539e-13, 1.825866e-13, 
    1.811974e-13, 1.824073e-13, 1.812158e-13, 1.812081e-13, 1.811842e-13, 
    1.811231e-13, 1.810358e-13, 1.808945e-13, 1.826416e-13, 1.826635e-13, 
    1.826235e-13, 1.825621e-13, 1.824983e-13, 1.824021e-13, 1.811694e-13, 
    1.811782e-13, 1.811971e-13, 1.812083e-13, 1.811808e-13, 1.812105e-13, 
    1.82599e-13, 1.824409e-13, 1.826714e-13, 1.82612e-13, 1.825659e-13, 
    1.825867e-13, 1.824698e-13, 1.824388e-13, 1.812025e-13, 1.811774e-13, 
    1.811412e-13, 1.81214e-13, 1.807575e-13, 1.809677e-13, 1.826708e-13, 
    1.826417e-13, 1.825237e-13, 1.825832e-13, 1.811676e-13, 1.811902e-13, 
    1.812038e-13, 1.812145e-13, 1.812152e-13, 1.812175e-13, 1.812123e-13, 
    1.812175e-13, 1.824019e-13, 1.811993e-13, 1.825386e-13, 1.824895e-13, 
    1.825126e-13, 1.825369e-13, 1.824586e-13, 1.811814e-13, 1.811822e-13, 
    1.811939e-13, 1.812142e-13, 1.81168e-13, 1.811245e-13, 1.812169e-13, 
    1.826076e-13, 1.82541e-13, 1.825308e-13, 1.825581e-13, 1.811882e-13, 
    1.824303e-13, 1.812175e-13, 1.812109e-13, 1.812168e-13, 1.81217e-13, 
    1.812165e-13, 1.812066e-13, 1.811954e-13, 1.824266e-13, 1.825009e-13, 
    1.825542e-13, 1.825423e-13, 1.824822e-13, 1.811838e-13, 1.812153e-13, 
    1.812114e-13, 1.812173e-13, 1.824108e-13, 1.812001e-13, 1.811872e-13, 
    1.812136e-13, 1.824658e-13, 1.812075e-13, 1.825078e-13, 1.824901e-13, 
    1.824319e-13, 1.81202e-13, 1.812089e-13, 1.812141e-13, 1.812112e-13, 
    1.811851e-13, 1.81179e-13, 1.824334e-13, 1.8245e-13, 1.82494e-13, 
    1.825282e-13, 1.82497e-13, 1.824625e-13, 1.811851e-13, 1.812127e-13, 
    1.812151e-13, 1.812111e-13, 1.811657e-13, 1.812059e-13, 1.811234e-13, 
    1.811986e-13, 1.810297e-13, 1.812099e-13, 1.812e-13, 1.824292e-13, 
    1.811692e-13, 1.811966e-13, 1.812167e-13, 1.812136e-13, 1.812154e-13, 
    1.811787e-13, 1.8248e-13, 1.825058e-13, 1.825511e-13, 1.825047e-13, 
    1.825086e-13, 1.82461e-13, 1.824767e-13, 1.811865e-13, 1.824209e-13, 
    1.812165e-13, 1.812155e-13, 1.811374e-13, 1.810303e-13, 1.808715e-13, 
    1.807845e-13, 1.80756e-13, 1.807437e-13 ;

 FCH4TOCO2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4_DFSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCOV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGEV =
  7.566927, 7.584713, 7.581267, 7.59555, 7.587664, 7.596979, 7.570558, 
    7.585398, 7.575937, 7.568562, 7.623105, 7.59619, 7.651288, 7.634079, 
    7.679165, 7.648578, 7.684998, 7.678385, 7.698424, 7.692685, 7.718223, 
    7.701074, 7.73156, 7.714154, 7.716856, 7.7005, 7.601656, 7.619739, 
    7.600573, 7.603154, 7.602008, 7.587809, 7.580578, 7.565606, 7.568334, 
    7.579351, 7.604316, 7.595897, 7.617222, 7.616742, 7.640441, 7.629751, 
    7.671416, 7.658321, 7.692925, 7.684648, 7.692527, 7.690145, 7.692558, 
    7.680423, 7.685618, 7.674962, 7.631743, 7.643904, 7.607615, 7.585694, 
    7.571198, 7.560875, 7.562334, 7.565104, 7.579414, 7.5929, 7.603112, 
    7.609937, 7.616672, 7.636908, 7.647741, 7.673686, 7.669359, 7.676723, 
    7.683826, 7.695698, 7.69375, 7.698971, 7.676562, 7.691436, 7.665132, 
    7.673591, 7.618323, 7.598176, 7.589461, 7.581923, 7.563452, 7.576197, 
    7.571168, 7.583172, 7.590768, 7.587023, 7.610124, 7.60114, 7.648383, 
    7.628031, 7.682998, 7.670251, 7.686062, 7.678, 7.691801, 7.67938, 
    7.700929, 7.705603, 7.702404, 7.714754, 7.678688, 7.69251, 7.586909, 
    7.58752, 7.590383, 7.577778, 7.577018, 7.565522, 7.575768, 7.580116, 
    7.59122, 7.597718, 7.603909, 7.617529, 7.632702, 7.653987, 7.671075, 
    7.681361, 7.675065, 7.680622, 7.674403, 7.671497, 7.70384, 7.685656, 
    7.712976, 7.71147, 7.699088, 7.71164, 7.587952, 7.58443, 7.572147, 
    7.581759, 7.564273, 7.574037, 7.579638, 7.601289, 7.606076, 7.61046, 
    7.61916, 7.630297, 7.649838, 7.668635, 7.684247, 7.683107, 7.683506, 
    7.686978, 7.678356, 7.688396, 7.690063, 7.685675, 7.711267, 7.703955, 
    7.711438, 7.706681, 7.58558, 7.591502, 7.588305, 7.594299, 7.590068, 
    7.608838, 7.614468, 7.640856, 7.630067, 7.647288, 7.631831, 7.634559, 
    7.647774, 7.632678, 7.667659, 7.643307, 7.687113, 7.662678, 7.688531, 
    7.68418, 7.691403, 7.697855, 7.706007, 7.721005, 7.717538, 7.730117, 
    7.600309, 7.607944, 7.607305, 7.615321, 7.621238, 7.634107, 7.654721, 
    7.646979, 7.661232, 7.664083, 7.642449, 7.655697, 7.61308, 7.61993, 
    7.615877, 7.600891, 7.648716, 7.62415, 7.671323, 7.656249, 7.69693, 
    7.67752, 7.715622, 7.731843, 7.74728, 7.765149, 7.612148, 7.606955, 
    7.616283, 7.62912, 7.641131, 7.657054, 7.658703, 7.661677, 7.671184, 
    7.677691, 7.662586, 7.679326, 7.62145, 7.650866, 7.604961, 7.61874, 
    7.628378, 7.624184, 7.646102, 7.651258, 7.673974, 7.661398, 7.727809, 
    7.69917, 7.778879, 7.75655, 7.605133, 7.612146, 7.636497, 7.624916, 
    7.658136, 7.668059, 7.674739, 7.683225, 7.684167, 7.689203, 7.680948, 
    7.68889, 7.657088, 7.672264, 7.633753, 7.642674, 7.638581, 7.634068, 
    7.647995, 7.662787, 7.663157, 7.669649, 7.682917, 7.658271, 7.731408, 
    7.687192, 7.619789, 7.633216, 7.635201, 7.629985, 7.665484, 7.652609, 
    7.689087, 7.679703, 7.695096, 7.68744, 7.686312, 7.676498, 7.670378, 
    7.653189, 7.640656, 7.630748, 7.633056, 7.643942, 7.663705, 7.684228, 
    7.680106, 7.693926, 7.655723, 7.672718, 7.665051, 7.682237, 7.646761, 
    7.677061, 7.639453, 7.642605, 7.652354, 7.673717, 7.67814, 7.682768, 
    7.679924, 7.664217, 7.661958, 7.65213, 7.649391, 7.641922, 7.635715, 
    7.641373, 7.647305, 7.664246, 7.681261, 7.697938, 7.702043, 7.721412, 
    7.705568, 7.731643, 7.709358, 7.748007, 7.678796, 7.708815, 7.652816, 
    7.658661, 7.670937, 7.695226, 7.682165, 7.697467, 7.661874, 7.64429, 
    7.63981, 7.631341, 7.640004, 7.639301, 7.647589, 7.644929, 7.664809, 
    7.65413, 7.686269, 7.69736, 7.728778, 7.748028, 7.767729, 7.776404, 
    7.77905, 7.780153 ;

 FGR =
  -370.322, -370.9913, -370.8614, -371.4004, -371.102, -371.4544, -370.4581, 
    -371.0174, -370.6606, -370.3829, -372.4434, -371.4245, -373.5011, 
    -372.8538, -374.4933, -373.3999, -374.7117, -374.4631, -375.2138, 
    -374.9988, -375.9571, -375.3131, -376.4557, -375.8038, -375.9054, 
    -375.2917, -371.6308, -372.3167, -371.5899, -371.6878, -371.6441, 
    -371.1078, -370.8364, -370.2716, -370.3743, -370.7896, -371.7318, 
    -371.4129, -372.2189, -372.2007, -373.0928, -372.6908, -374.2018, 
    -373.7639, -375.0078, -374.6977, -374.993, -374.9036, -374.9942, 
    -374.5396, -374.7343, -374.3346, -372.7659, -373.2232, -371.8563, 
    -371.0295, -370.4825, -370.0935, -370.1485, -370.2531, -370.792, 
    -371.2995, -371.6855, -371.9436, -372.1981, -372.9618, -373.368, 
    -374.2874, -374.1244, -374.4012, -374.6669, -375.1119, -375.0388, 
    -375.2347, -374.3946, -374.9526, -374.0194, -374.2832, -372.2635, 
    -371.4991, -371.171, -370.8862, -370.1907, -370.6708, -370.4814, 
    -370.9327, -371.2189, -371.0776, -371.9507, -371.6111, -373.392, 
    -372.6266, -374.636, -374.158, -374.7506, -374.4484, -374.9661, 
    -374.5002, -375.3079, -375.4834, -375.3634, -375.8256, -374.4742, 
    -374.9927, -371.0735, -371.0965, -371.2042, -370.7304, -370.7016, 
    -370.2686, -370.6542, -370.8182, -371.2358, -371.4818, -371.7159, 
    -372.2308, -372.8024, -373.602, -374.1889, -374.5743, -374.3382, 
    -374.5467, -374.3135, -374.2044, -375.4174, -374.7359, -375.7591, 
    -375.7026, -375.2392, -375.709, -371.1127, -370.98, -370.518, -370.8796, 
    -370.2215, -370.5893, -370.8006, -371.6174, -371.7976, -371.9636, 
    -372.292, -372.7113, -373.4461, -374.0977, -374.6825, -374.6397, 
    -374.6548, -374.7851, -374.4619, -374.8382, -374.901, -374.7362, 
    -375.695, -375.4211, -375.7014, -375.5232, -371.0233, -371.2466, 
    -371.1259, -371.3526, -371.1927, -371.903, -372.116, -373.1092, 
    -372.7029, -373.3505, -372.769, -372.8718, -373.3701, -372.8006, 
    -374.0618, -373.2017, -374.7902, -373.9294, -374.8433, -374.68, 
    -374.9507, -375.1928, -375.498, -376.0604, -375.9303, -376.4012, 
    -371.5797, -371.8688, -371.844, -372.1472, -372.3705, -372.8544, 
    -373.6291, -373.3382, -373.8731, -373.9803, -373.1678, -373.666, 
    -372.0629, -372.3221, -372.1684, -371.6021, -373.4043, -372.481, 
    -374.1983, -373.6863, -375.1582, -374.4313, -375.8585, -376.4672, 
    -377.0433, -377.7131, -372.0274, -371.8308, -372.1834, -372.6678, 
    -373.1187, -373.7167, -373.7782, -373.8901, -374.1927, -374.4368, 
    -373.9248, -374.498, -372.3807, -373.4847, -371.7559, -372.2774, 
    -372.6396, -372.4815, -373.3051, -373.4987, -374.2981, -373.8793, 
    -376.3164, -375.243, -378.2255, -377.3912, -371.762, -372.027, -372.9449, 
    -372.509, -373.757, -374.0758, -374.326, -374.6447, -374.6796, -374.8686, 
    -374.5589, -374.8566, -373.718, -374.2334, -372.8409, -373.1766, 
    -373.0224, -372.8528, -373.3762, -373.9325, -373.9455, -374.1357, 
    -374.6365, -373.762, -376.4531, -374.7963, -372.3156, -372.8221, 
    -372.8957, -372.6993, -374.033, -373.5497, -374.8641, -374.5122, 
    -375.0891, -374.8023, -374.7601, -374.3921, -374.1627, -373.5717, 
    -373.1009, -372.728, -372.8148, -373.2245, -373.9668, -374.6823, 
    -374.528, -375.0453, -373.6665, -374.2509, -374.0172, -374.6074, 
    -373.3302, -374.4163, -373.0552, -373.1737, -373.5402, -374.289, 
    -374.4536, -374.6276, -374.5205, -373.9859, -373.9007, -373.5315, 
    -373.4291, -373.148, -372.9147, -373.1276, -373.3509, -373.9865, 
    -374.5712, -375.1961, -375.3495, -376.0773, -375.4833, -376.4621, 
    -375.6278, -377.0733, -374.4802, -375.6053, -373.5572, -373.7766, 
    -374.1845, -375.0954, -374.6047, -375.1791, -373.8975, -373.2381, 
    -373.0687, -372.7505, -373.076, -373.0495, -373.3609, -373.2609, 
    -374.0076, -373.6065, -374.7588, -375.1748, -376.3514, -377.0724, 
    -377.8082, -378.1325, -378.2314, -378.2726 ;

 FGR12 =
  -167.3656, -167.4189, -167.4086, -167.4514, -167.4278, -167.4557, 
    -167.3765, -167.4209, -167.3926, -167.3706, -167.5341, -167.4534, 
    -167.6177, -167.567, -167.6965, -167.6097, -167.714, -167.6943, 
    -167.7543, -167.7371, -167.8138, -167.7623, -167.8542, -167.8016, 
    -167.8097, -167.7606, -167.4699, -167.5241, -167.4666, -167.4744, 
    -167.471, -167.4282, -167.4064, -167.3618, -167.3699, -167.4028, 
    -167.4779, -167.4526, -167.517, -167.5155, -167.5858, -167.5542, 
    -167.6735, -167.6386, -167.7378, -167.713, -167.7366, -167.7295, 
    -167.7367, -167.7004, -167.7159, -167.6841, -167.56, -167.5959, 
    -167.4879, -167.4217, -167.3784, -167.3476, -167.3519, -167.3602, 
    -167.403, -167.4436, -167.4743, -167.4949, -167.5153, -167.5751, 
    -167.6072, -167.6802, -167.6674, -167.6893, -167.7106, -167.7461, 
    -167.7403, -167.7559, -167.6889, -167.7333, -167.6589, -167.68, 
    -167.5199, -167.4595, -167.433, -167.4105, -167.3553, -167.3933, 
    -167.3783, -167.4143, -167.4371, -167.4259, -167.4955, -167.4684, 
    -167.6091, -167.549, -167.7081, -167.6701, -167.7173, -167.6932, 
    -167.7344, -167.6973, -167.7619, -167.7759, -167.7663, -167.8035, 
    -167.6953, -167.7365, -167.4256, -167.4274, -167.436, -167.3981, 
    -167.3958, -167.3615, -167.3921, -167.4051, -167.4386, -167.4581, 
    -167.4767, -167.5179, -167.5628, -167.6257, -167.6725, -167.7032, 
    -167.6844, -167.701, -167.6825, -167.6738, -167.7705, -167.716, 
    -167.7981, -167.7936, -167.7563, -167.7941, -167.4287, -167.4181, 
    -167.3813, -167.4101, -167.3578, -167.3869, -167.4036, -167.4687, 
    -167.4833, -167.4965, -167.5227, -167.5558, -167.6135, -167.6652, 
    -167.7119, -167.7085, -167.7097, -167.72, -167.6943, -167.7242, 
    -167.7292, -167.7161, -167.793, -167.771, -167.7935, -167.7792, 
    -167.4216, -167.4394, -167.4298, -167.4478, -167.435, -167.4915, 
    -167.5085, -167.5869, -167.5551, -167.6059, -167.5603, -167.5684, 
    -167.6072, -167.5629, -167.6622, -167.5941, -167.7204, -167.6514, 
    -167.7247, -167.7117, -167.7333, -167.7526, -167.7771, -167.8223, 
    -167.8119, -167.8499, -167.4659, -167.4888, -167.487, -167.5112, 
    -167.5289, -167.5671, -167.6279, -167.6051, -167.6473, -167.6557, 
    -167.5918, -167.6308, -167.5044, -167.5249, -167.5129, -167.4676, 
    -167.6101, -167.5375, -167.6732, -167.6325, -167.7498, -167.6917, 
    -167.8061, -167.855, -167.9021, -167.9565, -167.5016, -167.4859, 
    -167.5141, -167.5522, -167.5878, -167.6348, -167.6398, -167.6486, 
    -167.6729, -167.6923, -167.6512, -167.6971, -167.5293, -167.6165, 
    -167.4799, -167.5213, -167.55, -167.5376, -167.6026, -167.6178, 
    -167.6811, -167.6478, -167.8427, -167.7565, -167.9987, -167.9303, 
    -167.4805, -167.5016, -167.5741, -167.5398, -167.6381, -167.6635, 
    -167.6835, -167.7088, -167.7116, -167.7267, -167.702, -167.7257, 
    -167.6349, -167.6761, -167.5661, -167.5924, -167.5803, -167.567, 
    -167.6081, -167.6518, -167.653, -167.6682, -167.7075, -167.6385, 
    -167.8534, -167.7204, -167.5246, -167.5643, -167.5703, -167.5549, 
    -167.6599, -167.6217, -167.7263, -167.6983, -167.7443, -167.7214, 
    -167.718, -167.6887, -167.6704, -167.6234, -167.5864, -167.5572, 
    -167.564, -167.5961, -167.6546, -167.7117, -167.6994, -167.7408, 
    -167.631, -167.6774, -167.6586, -167.7058, -167.6045, -167.69, -167.5829, 
    -167.5922, -167.621, -167.6803, -167.6936, -167.7074, -167.6989, 
    -167.6561, -167.6494, -167.6203, -167.6122, -167.5902, -167.5719, 
    -167.5885, -167.606, -167.6562, -167.7029, -167.7528, -167.7652, 
    -167.8233, -167.7757, -167.8541, -167.7868, -167.904, -167.6954, 
    -167.7853, -167.6224, -167.6396, -167.672, -167.7446, -167.7056, 
    -167.7513, -167.6492, -167.5971, -167.5839, -167.5589, -167.5845, 
    -167.5824, -167.6069, -167.5991, -167.6579, -167.6262, -167.7179, 
    -167.7511, -167.8458, -167.9042, -167.9645, -167.9911, -167.9993, 
    -168.0027 ;

 FGR_R =
  -370.322, -370.9913, -370.8614, -371.4004, -371.102, -371.4544, -370.4581, 
    -371.0174, -370.6606, -370.3829, -372.4434, -371.4245, -373.5011, 
    -372.8538, -374.4933, -373.3999, -374.7117, -374.4631, -375.2138, 
    -374.9988, -375.9571, -375.3131, -376.4557, -375.8038, -375.9054, 
    -375.2917, -371.6308, -372.3167, -371.5899, -371.6878, -371.6441, 
    -371.1078, -370.8364, -370.2716, -370.3743, -370.7896, -371.7318, 
    -371.4129, -372.2189, -372.2007, -373.0928, -372.6908, -374.2018, 
    -373.7639, -375.0078, -374.6977, -374.993, -374.9036, -374.9942, 
    -374.5396, -374.7343, -374.3346, -372.7659, -373.2232, -371.8563, 
    -371.0295, -370.4825, -370.0935, -370.1485, -370.2531, -370.792, 
    -371.2995, -371.6855, -371.9436, -372.1981, -372.9618, -373.368, 
    -374.2874, -374.1244, -374.4012, -374.6669, -375.1119, -375.0388, 
    -375.2347, -374.3946, -374.9526, -374.0194, -374.2832, -372.2635, 
    -371.4991, -371.171, -370.8862, -370.1907, -370.6708, -370.4814, 
    -370.9327, -371.2189, -371.0776, -371.9507, -371.6111, -373.392, 
    -372.6266, -374.636, -374.158, -374.7506, -374.4484, -374.9661, 
    -374.5002, -375.3079, -375.4834, -375.3634, -375.8256, -374.4742, 
    -374.9927, -371.0735, -371.0965, -371.2042, -370.7304, -370.7016, 
    -370.2686, -370.6542, -370.8182, -371.2358, -371.4818, -371.7159, 
    -372.2308, -372.8024, -373.602, -374.1889, -374.5743, -374.3382, 
    -374.5467, -374.3135, -374.2044, -375.4174, -374.7359, -375.7591, 
    -375.7026, -375.2392, -375.709, -371.1127, -370.98, -370.518, -370.8796, 
    -370.2215, -370.5893, -370.8006, -371.6174, -371.7976, -371.9636, 
    -372.292, -372.7113, -373.4461, -374.0977, -374.6825, -374.6397, 
    -374.6548, -374.7851, -374.4619, -374.8382, -374.901, -374.7362, 
    -375.695, -375.4211, -375.7014, -375.5232, -371.0233, -371.2466, 
    -371.1259, -371.3526, -371.1927, -371.903, -372.116, -373.1092, 
    -372.7029, -373.3505, -372.769, -372.8718, -373.3701, -372.8006, 
    -374.0618, -373.2017, -374.7902, -373.9294, -374.8433, -374.68, 
    -374.9507, -375.1928, -375.498, -376.0604, -375.9303, -376.4012, 
    -371.5797, -371.8688, -371.844, -372.1472, -372.3705, -372.8544, 
    -373.6291, -373.3382, -373.8731, -373.9803, -373.1678, -373.666, 
    -372.0629, -372.3221, -372.1684, -371.6021, -373.4043, -372.481, 
    -374.1983, -373.6863, -375.1582, -374.4313, -375.8585, -376.4672, 
    -377.0433, -377.7131, -372.0274, -371.8308, -372.1834, -372.6678, 
    -373.1187, -373.7167, -373.7782, -373.8901, -374.1927, -374.4368, 
    -373.9248, -374.498, -372.3807, -373.4847, -371.7559, -372.2774, 
    -372.6396, -372.4815, -373.3051, -373.4987, -374.2981, -373.8793, 
    -376.3164, -375.243, -378.2255, -377.3912, -371.762, -372.027, -372.9449, 
    -372.509, -373.757, -374.0758, -374.326, -374.6447, -374.6796, -374.8686, 
    -374.5589, -374.8566, -373.718, -374.2334, -372.8409, -373.1766, 
    -373.0224, -372.8528, -373.3762, -373.9325, -373.9455, -374.1357, 
    -374.6365, -373.762, -376.4531, -374.7963, -372.3156, -372.8221, 
    -372.8957, -372.6993, -374.033, -373.5497, -374.8641, -374.5122, 
    -375.0891, -374.8023, -374.7601, -374.3921, -374.1627, -373.5717, 
    -373.1009, -372.728, -372.8148, -373.2245, -373.9668, -374.6823, 
    -374.528, -375.0453, -373.6665, -374.2509, -374.0172, -374.6074, 
    -373.3302, -374.4163, -373.0552, -373.1737, -373.5402, -374.289, 
    -374.4536, -374.6276, -374.5205, -373.9859, -373.9007, -373.5315, 
    -373.4291, -373.148, -372.9147, -373.1276, -373.3509, -373.9865, 
    -374.5712, -375.1961, -375.3495, -376.0773, -375.4833, -376.4621, 
    -375.6278, -377.0733, -374.4802, -375.6053, -373.5572, -373.7766, 
    -374.1845, -375.0954, -374.6047, -375.1791, -373.8975, -373.2381, 
    -373.0687, -372.7505, -373.076, -373.0495, -373.3609, -373.2609, 
    -374.0076, -373.6065, -374.7588, -375.1748, -376.3514, -377.0724, 
    -377.8082, -378.1325, -378.2314, -378.2726 ;

 FGR_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FIRA =
  77.93616, 77.98288, 77.97382, 78.01147, 77.99061, 78.01526, 77.94567, 
    77.9847, 77.95981, 77.94042, 78.08457, 78.01317, 78.15942, 78.11363, 
    78.22837, 78.15224, 78.24383, 78.22625, 78.27937, 78.26416, 78.33192, 
    78.2864, 78.36719, 78.3211, 78.32827, 78.28488, 78.02761, 78.07563, 
    78.02474, 78.03159, 78.02854, 77.991, 77.97207, 77.93265, 77.93982, 
    77.9688, 78.03468, 78.01236, 78.06877, 78.0675, 78.13054, 78.1021, 
    78.20776, 78.17806, 78.2648, 78.24286, 78.26375, 78.25743, 78.26383, 
    78.23166, 78.24545, 78.21716, 78.10741, 78.13976, 78.04339, 77.98554, 
    77.94737, 77.92022, 77.92406, 77.93136, 77.96897, 78.00442, 78.03144, 
    78.04951, 78.06731, 78.12125, 78.14999, 78.21381, 78.20229, 78.22186, 
    78.24068, 78.27216, 78.26699, 78.28085, 78.22141, 78.26088, 78.19616, 
    78.21352, 78.07188, 78.01839, 77.99541, 77.97555, 77.927, 77.96052, 
    77.9473, 77.9788, 77.99878, 77.98891, 78.05, 78.02624, 78.1517, 78.09756, 
    78.23849, 78.20466, 78.2466, 78.22521, 78.26184, 78.22888, 78.28603, 
    78.29843, 78.28995, 78.32265, 78.22704, 78.26373, 77.98862, 77.99023, 
    77.99775, 77.96468, 77.96267, 77.93244, 77.95936, 77.9708, 77.99996, 
    78.01718, 78.03357, 78.06961, 78.10999, 78.16657, 78.20685, 78.23413, 
    78.21742, 78.23217, 78.21567, 78.20795, 78.29376, 78.24555, 78.31795, 
    78.31395, 78.28117, 78.3144, 77.99136, 77.9821, 77.94985, 77.97509, 
    77.92915, 77.95483, 77.96957, 78.02666, 78.03929, 78.0509, 78.07394, 
    78.10356, 78.15553, 78.20039, 78.24178, 78.23876, 78.23982, 78.24904, 
    78.22617, 78.2528, 78.25724, 78.24558, 78.31341, 78.29404, 78.31387, 
    78.30125, 77.98512, 78.00072, 77.99228, 78.00814, 77.99694, 78.04666, 
    78.06156, 78.13168, 78.10296, 78.14876, 78.10764, 78.11491, 78.15013, 
    78.10988, 78.19783, 78.13822, 78.2494, 78.18974, 78.25316, 78.24161, 
    78.26076, 78.27789, 78.29948, 78.33923, 78.33004, 78.36334, 78.02403, 
    78.04427, 78.04254, 78.06375, 78.07947, 78.11368, 78.16851, 78.1479, 
    78.1858, 78.19338, 78.13585, 78.17112, 78.05785, 78.07604, 78.06524, 
    78.0256, 78.15257, 78.08725, 78.20751, 78.17256, 78.27544, 78.22399, 
    78.32497, 78.36799, 78.40874, 78.45605, 78.05537, 78.04161, 78.06629, 
    78.10047, 78.13237, 78.17471, 78.17908, 78.187, 78.20712, 78.2244, 
    78.18945, 78.22873, 78.08015, 78.15827, 78.03636, 78.07288, 78.09848, 
    78.0873, 78.14555, 78.15928, 78.21456, 78.18623, 78.35732, 78.28142, 
    78.49226, 78.4333, 78.0368, 78.05534, 78.12007, 78.08924, 78.17757, 
    78.19884, 78.21655, 78.23911, 78.24158, 78.25494, 78.23303, 78.2541, 
    78.1748, 78.21, 78.11273, 78.13647, 78.12556, 78.11357, 78.1506, 
    78.18999, 78.19092, 78.20308, 78.23846, 78.17793, 78.36695, 78.24978, 
    78.0756, 78.11137, 78.1166, 78.10271, 78.19711, 78.16289, 78.25463, 
    78.22974, 78.27055, 78.25026, 78.24727, 78.22123, 78.20499, 78.16444, 
    78.13111, 78.10474, 78.11088, 78.13985, 78.19241, 78.24176, 78.23084, 
    78.26746, 78.17116, 78.21123, 78.19599, 78.23647, 78.14733, 78.22289, 
    78.12788, 78.13627, 78.16221, 78.21391, 78.22559, 78.23789, 78.23032, 
    78.19377, 78.18774, 78.1616, 78.15434, 78.13445, 78.11795, 78.133, 
    78.1488, 78.19382, 78.23389, 78.27811, 78.28897, 78.34041, 78.29841, 
    78.36758, 78.30859, 78.41081, 78.22743, 78.30703, 78.16341, 78.17896, 
    78.20652, 78.27097, 78.23627, 78.2769, 78.18752, 78.1408, 78.12884, 
    78.10632, 78.12935, 78.12748, 78.14951, 78.14243, 78.19532, 78.16692, 
    78.24717, 78.2766, 78.35982, 78.41077, 78.46279, 78.4857, 78.49268, 
    78.4956 ;

 FIRA_R =
  77.93616, 77.98288, 77.97382, 78.01147, 77.99061, 78.01526, 77.94567, 
    77.9847, 77.95981, 77.94042, 78.08457, 78.01317, 78.15942, 78.11363, 
    78.22837, 78.15224, 78.24383, 78.22625, 78.27937, 78.26416, 78.33192, 
    78.2864, 78.36719, 78.3211, 78.32827, 78.28488, 78.02761, 78.07563, 
    78.02474, 78.03159, 78.02854, 77.991, 77.97207, 77.93265, 77.93982, 
    77.9688, 78.03468, 78.01236, 78.06877, 78.0675, 78.13054, 78.1021, 
    78.20776, 78.17806, 78.2648, 78.24286, 78.26375, 78.25743, 78.26383, 
    78.23166, 78.24545, 78.21716, 78.10741, 78.13976, 78.04339, 77.98554, 
    77.94737, 77.92022, 77.92406, 77.93136, 77.96897, 78.00442, 78.03144, 
    78.04951, 78.06731, 78.12125, 78.14999, 78.21381, 78.20229, 78.22186, 
    78.24068, 78.27216, 78.26699, 78.28085, 78.22141, 78.26088, 78.19616, 
    78.21352, 78.07188, 78.01839, 77.99541, 77.97555, 77.927, 77.96052, 
    77.9473, 77.9788, 77.99878, 77.98891, 78.05, 78.02624, 78.1517, 78.09756, 
    78.23849, 78.20466, 78.2466, 78.22521, 78.26184, 78.22888, 78.28603, 
    78.29843, 78.28995, 78.32265, 78.22704, 78.26373, 77.98862, 77.99023, 
    77.99775, 77.96468, 77.96267, 77.93244, 77.95936, 77.9708, 77.99996, 
    78.01718, 78.03357, 78.06961, 78.10999, 78.16657, 78.20685, 78.23413, 
    78.21742, 78.23217, 78.21567, 78.20795, 78.29376, 78.24555, 78.31795, 
    78.31395, 78.28117, 78.3144, 77.99136, 77.9821, 77.94985, 77.97509, 
    77.92915, 77.95483, 77.96957, 78.02666, 78.03929, 78.0509, 78.07394, 
    78.10356, 78.15553, 78.20039, 78.24178, 78.23876, 78.23982, 78.24904, 
    78.22617, 78.2528, 78.25724, 78.24558, 78.31341, 78.29404, 78.31387, 
    78.30125, 77.98512, 78.00072, 77.99228, 78.00814, 77.99694, 78.04666, 
    78.06156, 78.13168, 78.10296, 78.14876, 78.10764, 78.11491, 78.15013, 
    78.10988, 78.19783, 78.13822, 78.2494, 78.18974, 78.25316, 78.24161, 
    78.26076, 78.27789, 78.29948, 78.33923, 78.33004, 78.36334, 78.02403, 
    78.04427, 78.04254, 78.06375, 78.07947, 78.11368, 78.16851, 78.1479, 
    78.1858, 78.19338, 78.13585, 78.17112, 78.05785, 78.07604, 78.06524, 
    78.0256, 78.15257, 78.08725, 78.20751, 78.17256, 78.27544, 78.22399, 
    78.32497, 78.36799, 78.40874, 78.45605, 78.05537, 78.04161, 78.06629, 
    78.10047, 78.13237, 78.17471, 78.17908, 78.187, 78.20712, 78.2244, 
    78.18945, 78.22873, 78.08015, 78.15827, 78.03636, 78.07288, 78.09848, 
    78.0873, 78.14555, 78.15928, 78.21456, 78.18623, 78.35732, 78.28142, 
    78.49226, 78.4333, 78.0368, 78.05534, 78.12007, 78.08924, 78.17757, 
    78.19884, 78.21655, 78.23911, 78.24158, 78.25494, 78.23303, 78.2541, 
    78.1748, 78.21, 78.11273, 78.13647, 78.12556, 78.11357, 78.1506, 
    78.18999, 78.19092, 78.20308, 78.23846, 78.17793, 78.36695, 78.24978, 
    78.0756, 78.11137, 78.1166, 78.10271, 78.19711, 78.16289, 78.25463, 
    78.22974, 78.27055, 78.25026, 78.24727, 78.22123, 78.20499, 78.16444, 
    78.13111, 78.10474, 78.11088, 78.13985, 78.19241, 78.24176, 78.23084, 
    78.26746, 78.17116, 78.21123, 78.19599, 78.23647, 78.14733, 78.22289, 
    78.12788, 78.13627, 78.16221, 78.21391, 78.22559, 78.23789, 78.23032, 
    78.19377, 78.18774, 78.1616, 78.15434, 78.13445, 78.11795, 78.133, 
    78.1488, 78.19382, 78.23389, 78.27811, 78.28897, 78.34041, 78.29841, 
    78.36758, 78.30859, 78.41081, 78.22743, 78.30703, 78.16341, 78.17896, 
    78.20652, 78.27097, 78.23627, 78.2769, 78.18752, 78.1408, 78.12884, 
    78.10632, 78.12935, 78.12748, 78.14951, 78.14243, 78.19532, 78.16692, 
    78.24717, 78.2766, 78.35982, 78.41077, 78.46279, 78.4857, 78.49268, 
    78.4956 ;

 FIRA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FIRE =
  266.8971, 266.9438, 266.9348, 266.9724, 266.9515, 266.9762, 266.9066, 
    266.9456, 266.9207, 266.9014, 267.0455, 266.9741, 267.1204, 267.0746, 
    267.1893, 267.1132, 267.2048, 267.1872, 267.2403, 267.2251, 267.2928, 
    267.2473, 267.3281, 267.282, 267.2892, 267.2458, 266.9886, 267.0366, 
    266.9857, 266.9925, 266.9895, 266.9519, 266.933, 266.8936, 266.9008, 
    266.9297, 266.9956, 266.9733, 267.0297, 267.0284, 267.0915, 267.063, 
    267.1687, 267.139, 267.2257, 267.2038, 267.2247, 267.2184, 267.2248, 
    267.1926, 267.2064, 267.1781, 267.0684, 267.1007, 267.0043, 266.9465, 
    266.9083, 266.8812, 266.885, 266.8923, 266.9299, 266.9654, 266.9924, 
    267.0104, 267.0283, 267.0822, 267.1109, 267.1747, 267.1632, 267.1828, 
    267.2016, 267.2331, 267.2279, 267.2418, 267.1823, 267.2218, 267.1571, 
    267.1745, 267.0328, 266.9793, 266.9564, 266.9365, 266.8879, 266.9214, 
    266.9082, 266.9397, 266.9597, 266.9499, 267.0109, 266.9872, 267.1126, 
    267.0585, 267.1994, 267.1656, 267.2076, 267.1862, 267.2228, 267.1898, 
    267.247, 267.2594, 267.2509, 267.2836, 267.188, 267.2247, 266.9496, 
    266.9512, 266.9587, 266.9256, 266.9236, 266.8934, 266.9203, 266.9317, 
    266.9609, 266.9781, 266.9945, 267.0305, 267.0709, 267.1275, 267.1678, 
    267.1951, 267.1783, 267.1931, 267.1766, 267.1689, 267.2547, 267.2065, 
    267.2789, 267.2749, 267.2421, 267.2753, 266.9523, 266.943, 266.9108, 
    266.936, 266.8901, 266.9158, 266.9305, 266.9876, 267.0002, 267.0118, 
    267.0349, 267.0645, 267.1165, 267.1613, 267.2027, 267.1997, 267.2008, 
    267.21, 267.1871, 267.2137, 267.2182, 267.2065, 267.2744, 267.255, 
    267.2748, 267.2622, 266.946, 266.9617, 266.9532, 266.9691, 266.9579, 
    267.0076, 267.0225, 267.0926, 267.0639, 267.1097, 267.0686, 267.0758, 
    267.1111, 267.0708, 267.1588, 267.0992, 267.2103, 267.1507, 267.2141, 
    267.2025, 267.2217, 267.2388, 267.2604, 267.3002, 267.291, 267.3243, 
    266.985, 267.0052, 267.0035, 267.0247, 267.0404, 267.0746, 267.1295, 
    267.1088, 267.1467, 267.1543, 267.0968, 267.132, 267.0188, 267.037, 
    267.0262, 266.9865, 267.1135, 267.0482, 267.1685, 267.1335, 267.2364, 
    267.1849, 267.2859, 267.3289, 267.3697, 267.417, 267.0163, 267.0026, 
    267.0272, 267.0614, 267.0933, 267.1357, 267.14, 267.1479, 267.1681, 
    267.1853, 267.1504, 267.1897, 267.0411, 267.1192, 266.9973, 267.0338, 
    267.0594, 267.0482, 267.1065, 267.1202, 267.1755, 267.1472, 267.3183, 
    267.2424, 267.4532, 267.3943, 266.9977, 267.0163, 267.081, 267.0502, 
    267.1385, 267.1598, 267.1775, 267.2, 267.2025, 267.2159, 267.194, 
    267.215, 267.1357, 267.1709, 267.0737, 267.0974, 267.0865, 267.0745, 
    267.1115, 267.1509, 267.1519, 267.164, 267.1994, 267.1389, 267.3279, 
    267.2107, 267.0365, 267.0723, 267.0775, 267.0637, 267.1581, 267.1238, 
    267.2156, 267.1907, 267.2315, 267.2112, 267.2082, 267.1822, 267.1659, 
    267.1254, 267.092, 267.0657, 267.0718, 267.1008, 267.1534, 267.2027, 
    267.1918, 267.2284, 267.1321, 267.1721, 267.1569, 267.1974, 267.1083, 
    267.1838, 267.0888, 267.0972, 267.1231, 267.1749, 267.1865, 267.1988, 
    267.1913, 267.1547, 267.1487, 267.1225, 267.1153, 267.0954, 267.0789, 
    267.0939, 267.1097, 267.1548, 267.1948, 267.239, 267.2499, 267.3013, 
    267.2593, 267.3285, 267.2695, 267.3718, 267.1884, 267.268, 267.1244, 
    267.1399, 267.1674, 267.2319, 267.1972, 267.2378, 267.1485, 267.1017, 
    267.0898, 267.0673, 267.0903, 267.0884, 267.1104, 267.1034, 267.1562, 
    267.1278, 267.2081, 267.2375, 267.3208, 267.3717, 267.4237, 267.4467, 
    267.4536, 267.4565 ;

 FIRE_R =
  266.8971, 266.9438, 266.9348, 266.9724, 266.9515, 266.9762, 266.9066, 
    266.9456, 266.9207, 266.9014, 267.0455, 266.9741, 267.1204, 267.0746, 
    267.1893, 267.1132, 267.2048, 267.1872, 267.2403, 267.2251, 267.2928, 
    267.2473, 267.3281, 267.282, 267.2892, 267.2458, 266.9886, 267.0366, 
    266.9857, 266.9925, 266.9895, 266.9519, 266.933, 266.8936, 266.9008, 
    266.9297, 266.9956, 266.9733, 267.0297, 267.0284, 267.0915, 267.063, 
    267.1687, 267.139, 267.2257, 267.2038, 267.2247, 267.2184, 267.2248, 
    267.1926, 267.2064, 267.1781, 267.0684, 267.1007, 267.0043, 266.9465, 
    266.9083, 266.8812, 266.885, 266.8923, 266.9299, 266.9654, 266.9924, 
    267.0104, 267.0283, 267.0822, 267.1109, 267.1747, 267.1632, 267.1828, 
    267.2016, 267.2331, 267.2279, 267.2418, 267.1823, 267.2218, 267.1571, 
    267.1745, 267.0328, 266.9793, 266.9564, 266.9365, 266.8879, 266.9214, 
    266.9082, 266.9397, 266.9597, 266.9499, 267.0109, 266.9872, 267.1126, 
    267.0585, 267.1994, 267.1656, 267.2076, 267.1862, 267.2228, 267.1898, 
    267.247, 267.2594, 267.2509, 267.2836, 267.188, 267.2247, 266.9496, 
    266.9512, 266.9587, 266.9256, 266.9236, 266.8934, 266.9203, 266.9317, 
    266.9609, 266.9781, 266.9945, 267.0305, 267.0709, 267.1275, 267.1678, 
    267.1951, 267.1783, 267.1931, 267.1766, 267.1689, 267.2547, 267.2065, 
    267.2789, 267.2749, 267.2421, 267.2753, 266.9523, 266.943, 266.9108, 
    266.936, 266.8901, 266.9158, 266.9305, 266.9876, 267.0002, 267.0118, 
    267.0349, 267.0645, 267.1165, 267.1613, 267.2027, 267.1997, 267.2008, 
    267.21, 267.1871, 267.2137, 267.2182, 267.2065, 267.2744, 267.255, 
    267.2748, 267.2622, 266.946, 266.9617, 266.9532, 266.9691, 266.9579, 
    267.0076, 267.0225, 267.0926, 267.0639, 267.1097, 267.0686, 267.0758, 
    267.1111, 267.0708, 267.1588, 267.0992, 267.2103, 267.1507, 267.2141, 
    267.2025, 267.2217, 267.2388, 267.2604, 267.3002, 267.291, 267.3243, 
    266.985, 267.0052, 267.0035, 267.0247, 267.0404, 267.0746, 267.1295, 
    267.1088, 267.1467, 267.1543, 267.0968, 267.132, 267.0188, 267.037, 
    267.0262, 266.9865, 267.1135, 267.0482, 267.1685, 267.1335, 267.2364, 
    267.1849, 267.2859, 267.3289, 267.3697, 267.417, 267.0163, 267.0026, 
    267.0272, 267.0614, 267.0933, 267.1357, 267.14, 267.1479, 267.1681, 
    267.1853, 267.1504, 267.1897, 267.0411, 267.1192, 266.9973, 267.0338, 
    267.0594, 267.0482, 267.1065, 267.1202, 267.1755, 267.1472, 267.3183, 
    267.2424, 267.4532, 267.3943, 266.9977, 267.0163, 267.081, 267.0502, 
    267.1385, 267.1598, 267.1775, 267.2, 267.2025, 267.2159, 267.194, 
    267.215, 267.1357, 267.1709, 267.0737, 267.0974, 267.0865, 267.0745, 
    267.1115, 267.1509, 267.1519, 267.164, 267.1994, 267.1389, 267.3279, 
    267.2107, 267.0365, 267.0723, 267.0775, 267.0637, 267.1581, 267.1238, 
    267.2156, 267.1907, 267.2315, 267.2112, 267.2082, 267.1822, 267.1659, 
    267.1254, 267.092, 267.0657, 267.0718, 267.1008, 267.1534, 267.2027, 
    267.1918, 267.2284, 267.1321, 267.1721, 267.1569, 267.1974, 267.1083, 
    267.1838, 267.0888, 267.0972, 267.1231, 267.1749, 267.1865, 267.1988, 
    267.1913, 267.1547, 267.1487, 267.1225, 267.1153, 267.0954, 267.0789, 
    267.0939, 267.1097, 267.1548, 267.1948, 267.239, 267.2499, 267.3013, 
    267.2593, 267.3285, 267.2695, 267.3718, 267.1884, 267.268, 267.1244, 
    267.1399, 267.1674, 267.2319, 267.1972, 267.2378, 267.1485, 267.1017, 
    267.0898, 267.0673, 267.0903, 267.0884, 267.1104, 267.1034, 267.1562, 
    267.1278, 267.2081, 267.2375, 267.3208, 267.3717, 267.4237, 267.4467, 
    267.4536, 267.4565 ;

 FIRE_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FLDS =
  188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609 ;

 FPG =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI_vr =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WJ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROST_TABLE =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 FSA =
  0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643 ;

 FSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSA_R =
  0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643 ;

 FSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSDS =
  1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658 ;

 FSDSND =
  0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004 ;

 FSDSNDLN =
  0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372 ;

 FSDSNI =
  0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284 ;

 FSDSVD =
  0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081 ;

 FSDSVDLN =
  0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678 ;

 FSDSVI =
  0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228 ;

 FSDSVILN =
  0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012 ;

 FSH =
  286.4722, 287.0759, 286.9588, 287.4449, 287.1758, 287.4937, 286.595, 
    287.0995, 286.7777, 286.5271, 288.3857, 287.4667, 289.3385, 288.7552, 
    290.2322, 289.2473, 290.429, 290.205, 290.8813, 290.6875, 291.551, 
    290.9707, 292.0001, 291.4128, 291.5044, 290.9514, 287.6527, 288.2714, 
    287.6158, 287.7041, 287.6647, 287.181, 286.9363, 286.4267, 286.5194, 
    286.894, 287.7439, 287.4561, 288.1831, 288.1667, 288.9706, 288.6083, 
    289.9695, 289.5752, 290.6956, 290.4164, 290.6824, 290.6018, 290.6834, 
    290.2739, 290.4493, 290.0892, 288.676, 289.0881, 287.8561, 287.1105, 
    286.617, 286.2661, 286.3157, 286.4101, 286.8962, 287.3539, 287.7021, 
    287.9348, 288.1643, 288.8527, 289.2186, 290.0468, 289.8999, 290.1493, 
    290.3886, 290.7895, 290.7236, 290.9001, 290.1432, 290.6459, 289.8053, 
    290.0429, 288.2235, 287.5339, 287.2381, 286.9812, 286.3538, 286.7869, 
    286.6161, 287.0231, 287.2812, 287.1537, 287.9412, 287.6349, 289.2402, 
    288.5506, 290.3607, 289.9301, 290.464, 290.1917, 290.6581, 290.2383, 
    290.966, 291.1242, 291.016, 291.4324, 290.215, 290.6821, 287.15, 
    287.1708, 287.268, 286.8406, 286.8147, 286.424, 286.7719, 286.9198, 
    287.2964, 287.5183, 287.7295, 288.1938, 288.709, 289.4293, 289.9579, 
    290.3052, 290.0924, 290.2802, 290.0702, 289.9719, 291.0647, 290.4507, 
    291.3725, 291.3216, 290.9042, 291.3274, 287.1855, 287.0657, 286.649, 
    286.9751, 286.3815, 286.7134, 286.904, 287.6407, 287.8032, 287.9529, 
    288.249, 288.6269, 289.2889, 289.8758, 290.4026, 290.3641, 290.3776, 
    290.4951, 290.2038, 290.5429, 290.5995, 290.451, 291.3148, 291.068, 
    291.3205, 291.1599, 287.1047, 287.3062, 287.1974, 287.4019, 287.2576, 
    287.8983, 288.0904, 288.9854, 288.6193, 289.2028, 288.6788, 288.7715, 
    289.2206, 288.7073, 289.8435, 289.0688, 290.4996, 289.7243, 290.5475, 
    290.4004, 290.6442, 290.8623, 291.1373, 291.644, 291.5267, 291.951, 
    287.6066, 287.8674, 287.845, 288.1184, 288.3198, 288.7558, 289.4538, 
    289.1916, 289.6736, 289.7702, 289.0382, 289.4871, 288.0424, 288.2762, 
    288.1376, 287.6268, 289.2513, 288.4193, 289.9664, 289.5053, 290.8311, 
    290.1764, 291.4621, 292.0106, 292.5294, 293.133, 288.0104, 287.8331, 
    288.1511, 288.5878, 288.9939, 289.5327, 289.5881, 289.6888, 289.9613, 
    290.1812, 289.7202, 290.2364, 288.3291, 289.3237, 287.7655, 288.2359, 
    288.5623, 288.4198, 289.1618, 289.3363, 290.0563, 289.6791, 291.8747, 
    290.9077, 293.5944, 292.8429, 287.771, 288.0101, 288.8374, 288.4445, 
    289.5689, 289.8561, 290.0814, 290.3686, 290.4, 290.5703, 290.2912, 
    290.5595, 289.5338, 289.998, 288.7436, 289.0461, 288.9072, 288.7543, 
    289.2259, 289.7271, 289.7387, 289.9101, 290.3614, 289.5735, 291.9979, 
    290.5053, 288.2703, 288.7267, 288.793, 288.6161, 289.8176, 289.3823, 
    290.5663, 290.2492, 290.769, 290.5106, 290.4725, 290.141, 289.9344, 
    289.402, 288.9779, 288.6418, 288.7201, 289.0892, 289.758, 290.4025, 
    290.2635, 290.7295, 289.4874, 290.0138, 289.8034, 290.335, 289.1845, 
    290.163, 288.9367, 289.0435, 289.3736, 290.0482, 290.1964, 290.3532, 
    290.2567, 289.7752, 289.6985, 289.3658, 289.2736, 289.0203, 288.8101, 
    289.0019, 289.2032, 289.7757, 290.3023, 290.8653, 291.0034, 291.6593, 
    291.1242, 292.0061, 291.2545, 292.5566, 290.2204, 291.2341, 289.3889, 
    289.5866, 289.9541, 290.7747, 290.3325, 290.85, 289.6955, 289.1015, 
    288.9488, 288.6621, 288.9554, 288.9316, 289.2121, 289.122, 289.7948, 
    289.4334, 290.4713, 290.8462, 291.9062, 292.5557, 293.2185, 293.5107, 
    293.5997, 293.6369 ;

 FSH_G =
  299.5754, 300.1801, 300.0627, 300.5497, 300.2801, 300.5985, 299.6984, 
    300.2037, 299.8814, 299.6304, 301.4919, 300.5715, 302.4464, 301.8622, 
    303.3415, 302.3551, 303.5386, 303.3143, 303.9916, 303.7976, 304.6624, 
    304.0812, 305.1123, 304.5241, 304.6158, 304.0619, 300.7578, 301.3775, 
    300.7209, 300.8093, 300.7698, 300.2853, 300.0402, 299.5298, 299.6227, 
    299.9979, 300.8491, 300.5609, 301.2891, 301.2727, 302.0779, 301.7151, 
    303.0785, 302.6835, 303.8057, 303.526, 303.7924, 303.7118, 303.7935, 
    303.3832, 303.559, 303.1983, 301.7828, 302.1956, 300.9615, 300.2147, 
    299.7204, 299.369, 299.4187, 299.5132, 300, 300.4586, 300.8073, 301.0404, 
    301.2703, 301.9597, 302.3262, 303.1558, 303.0086, 303.2584, 303.4982, 
    303.8997, 303.8337, 304.0105, 303.2524, 303.7559, 302.914, 303.1519, 
    301.3296, 300.6388, 300.3425, 300.0852, 299.4568, 299.8905, 299.7195, 
    300.1272, 300.3858, 300.2581, 301.0468, 300.7401, 302.3479, 301.6572, 
    303.4702, 303.0389, 303.5737, 303.3009, 303.7681, 303.3477, 304.0765, 
    304.235, 304.1266, 304.5438, 303.3243, 303.7921, 300.2543, 300.2751, 
    300.3725, 299.9444, 299.9184, 299.5271, 299.8756, 300.0237, 300.401, 
    300.6232, 300.8347, 301.2999, 301.8158, 302.5374, 303.0668, 303.4146, 
    303.2015, 303.3896, 303.1793, 303.0808, 304.1754, 303.5604, 304.4837, 
    304.4327, 304.0146, 304.4385, 300.2898, 300.1699, 299.7525, 300.0791, 
    299.4846, 299.817, 300.0078, 300.7458, 300.9086, 301.0585, 301.3551, 
    301.7336, 302.3967, 302.9846, 303.5122, 303.4736, 303.4872, 303.6048, 
    303.3131, 303.6527, 303.7094, 303.5607, 304.4259, 304.1787, 304.4317, 
    304.2708, 300.209, 300.4108, 300.3017, 300.5066, 300.3621, 301.0038, 
    301.1963, 302.0927, 301.726, 302.3105, 301.7856, 301.8784, 302.3282, 
    301.8142, 302.9521, 302.1762, 303.6094, 302.8328, 303.6573, 303.5099, 
    303.7542, 303.9727, 304.2481, 304.7556, 304.6382, 305.0631, 300.7116, 
    300.9729, 300.9505, 301.2243, 301.426, 301.8627, 302.5619, 302.2993, 
    302.782, 302.8788, 302.1456, 302.5952, 301.1482, 301.3823, 301.2435, 
    300.7319, 302.359, 301.5257, 303.0753, 302.6135, 303.9415, 303.2856, 
    304.5734, 305.1228, 305.6425, 306.2471, 301.1161, 300.9385, 301.2571, 
    301.6944, 302.1013, 302.6409, 302.6964, 302.7973, 303.0702, 303.2905, 
    302.8287, 303.3458, 301.4353, 302.4315, 300.8708, 301.342, 301.6689, 
    301.5262, 302.2694, 302.4442, 303.1653, 302.7876, 304.9867, 304.0181, 
    306.7093, 305.9565, 300.8763, 301.1158, 301.9444, 301.551, 302.6772, 
    302.9648, 303.1905, 303.4781, 303.5096, 303.6801, 303.4007, 303.6693, 
    302.642, 303.107, 301.8506, 302.1535, 302.0143, 301.8613, 302.3336, 
    302.8357, 302.8473, 303.0189, 303.4709, 302.6818, 305.1101, 303.615, 
    301.3764, 301.8336, 301.9, 301.7228, 302.9263, 302.4902, 303.6761, 
    303.3586, 303.8792, 303.6204, 303.5822, 303.2502, 303.0432, 302.51, 
    302.0852, 301.7486, 301.8269, 302.1967, 302.8666, 303.5121, 303.3729, 
    303.8396, 302.5955, 303.1227, 302.9121, 303.4445, 302.2921, 303.2722, 
    302.0439, 302.1509, 302.4816, 303.1572, 303.3057, 303.4627, 303.366, 
    302.8838, 302.8069, 302.4738, 302.3813, 302.1277, 301.9171, 302.1093, 
    302.3108, 302.8843, 303.4118, 303.9757, 304.114, 304.7709, 304.235, 
    305.1183, 304.3654, 305.6697, 303.3297, 304.3451, 302.4969, 302.6949, 
    303.0629, 303.8849, 303.442, 303.9604, 302.804, 302.209, 302.0561, 
    301.7689, 302.0627, 302.0388, 302.3198, 302.2296, 302.9034, 302.5414, 
    303.5811, 303.9565, 305.0182, 305.6689, 306.3328, 306.6255, 306.7146, 
    306.7519 ;

 FSH_NODYNLNDUSE =
  286.4722, 287.0759, 286.9588, 287.4449, 287.1758, 287.4937, 286.595, 
    287.0995, 286.7777, 286.5271, 288.3857, 287.4667, 289.3385, 288.7552, 
    290.2322, 289.2473, 290.429, 290.205, 290.8813, 290.6875, 291.551, 
    290.9707, 292.0001, 291.4128, 291.5044, 290.9514, 287.6527, 288.2714, 
    287.6158, 287.7041, 287.6647, 287.181, 286.9363, 286.4267, 286.5194, 
    286.894, 287.7439, 287.4561, 288.1831, 288.1667, 288.9706, 288.6083, 
    289.9695, 289.5752, 290.6956, 290.4164, 290.6824, 290.6018, 290.6834, 
    290.2739, 290.4493, 290.0892, 288.676, 289.0881, 287.8561, 287.1105, 
    286.617, 286.2661, 286.3157, 286.4101, 286.8962, 287.3539, 287.7021, 
    287.9348, 288.1643, 288.8527, 289.2186, 290.0468, 289.8999, 290.1493, 
    290.3886, 290.7895, 290.7236, 290.9001, 290.1432, 290.6459, 289.8053, 
    290.0429, 288.2235, 287.5339, 287.2381, 286.9812, 286.3538, 286.7869, 
    286.6161, 287.0231, 287.2812, 287.1537, 287.9412, 287.6349, 289.2402, 
    288.5506, 290.3607, 289.9301, 290.464, 290.1917, 290.6581, 290.2383, 
    290.966, 291.1242, 291.016, 291.4324, 290.215, 290.6821, 287.15, 
    287.1708, 287.268, 286.8406, 286.8147, 286.424, 286.7719, 286.9198, 
    287.2964, 287.5183, 287.7295, 288.1938, 288.709, 289.4293, 289.9579, 
    290.3052, 290.0924, 290.2802, 290.0702, 289.9719, 291.0647, 290.4507, 
    291.3725, 291.3216, 290.9042, 291.3274, 287.1855, 287.0657, 286.649, 
    286.9751, 286.3815, 286.7134, 286.904, 287.6407, 287.8032, 287.9529, 
    288.249, 288.6269, 289.2889, 289.8758, 290.4026, 290.3641, 290.3776, 
    290.4951, 290.2038, 290.5429, 290.5995, 290.451, 291.3148, 291.068, 
    291.3205, 291.1599, 287.1047, 287.3062, 287.1974, 287.4019, 287.2576, 
    287.8983, 288.0904, 288.9854, 288.6193, 289.2028, 288.6788, 288.7715, 
    289.2206, 288.7073, 289.8435, 289.0688, 290.4996, 289.7243, 290.5475, 
    290.4004, 290.6442, 290.8623, 291.1373, 291.644, 291.5267, 291.951, 
    287.6066, 287.8674, 287.845, 288.1184, 288.3198, 288.7558, 289.4538, 
    289.1916, 289.6736, 289.7702, 289.0382, 289.4871, 288.0424, 288.2762, 
    288.1376, 287.6268, 289.2513, 288.4193, 289.9664, 289.5053, 290.8311, 
    290.1764, 291.4621, 292.0106, 292.5294, 293.133, 288.0104, 287.8331, 
    288.1511, 288.5878, 288.9939, 289.5327, 289.5881, 289.6888, 289.9613, 
    290.1812, 289.7202, 290.2364, 288.3291, 289.3237, 287.7655, 288.2359, 
    288.5623, 288.4198, 289.1618, 289.3363, 290.0563, 289.6791, 291.8747, 
    290.9077, 293.5944, 292.8429, 287.771, 288.0101, 288.8374, 288.4445, 
    289.5689, 289.8561, 290.0814, 290.3686, 290.4, 290.5703, 290.2912, 
    290.5595, 289.5338, 289.998, 288.7436, 289.0461, 288.9072, 288.7543, 
    289.2259, 289.7271, 289.7387, 289.9101, 290.3614, 289.5735, 291.9979, 
    290.5053, 288.2703, 288.7267, 288.793, 288.6161, 289.8176, 289.3823, 
    290.5663, 290.2492, 290.769, 290.5106, 290.4725, 290.141, 289.9344, 
    289.402, 288.9779, 288.6418, 288.7201, 289.0892, 289.758, 290.4025, 
    290.2635, 290.7295, 289.4874, 290.0138, 289.8034, 290.335, 289.1845, 
    290.163, 288.9367, 289.0435, 289.3736, 290.0482, 290.1964, 290.3532, 
    290.2567, 289.7752, 289.6985, 289.3658, 289.2736, 289.0203, 288.8101, 
    289.0019, 289.2032, 289.7757, 290.3023, 290.8653, 291.0034, 291.6593, 
    291.1242, 292.0061, 291.2545, 292.5566, 290.2204, 291.2341, 289.3889, 
    289.5866, 289.9541, 290.7747, 290.3325, 290.85, 289.6955, 289.1015, 
    288.9488, 288.6621, 288.9554, 288.9316, 289.2121, 289.122, 289.7948, 
    289.4334, 290.4713, 290.8462, 291.9062, 292.5557, 293.2185, 293.5107, 
    293.5997, 293.6369 ;

 FSH_R =
  286.4722, 287.0759, 286.9588, 287.4449, 287.1758, 287.4937, 286.595, 
    287.0995, 286.7777, 286.5271, 288.3857, 287.4667, 289.3385, 288.7552, 
    290.2322, 289.2473, 290.429, 290.205, 290.8813, 290.6875, 291.551, 
    290.9707, 292.0001, 291.4128, 291.5044, 290.9514, 287.6527, 288.2714, 
    287.6158, 287.7041, 287.6647, 287.181, 286.9363, 286.4267, 286.5194, 
    286.894, 287.7439, 287.4561, 288.1831, 288.1667, 288.9706, 288.6083, 
    289.9695, 289.5752, 290.6956, 290.4164, 290.6824, 290.6018, 290.6834, 
    290.2739, 290.4493, 290.0892, 288.676, 289.0881, 287.8561, 287.1105, 
    286.617, 286.2661, 286.3157, 286.4101, 286.8962, 287.3539, 287.7021, 
    287.9348, 288.1643, 288.8527, 289.2186, 290.0468, 289.8999, 290.1493, 
    290.3886, 290.7895, 290.7236, 290.9001, 290.1432, 290.6459, 289.8053, 
    290.0429, 288.2235, 287.5339, 287.2381, 286.9812, 286.3538, 286.7869, 
    286.6161, 287.0231, 287.2812, 287.1537, 287.9412, 287.6349, 289.2402, 
    288.5506, 290.3607, 289.9301, 290.464, 290.1917, 290.6581, 290.2383, 
    290.966, 291.1242, 291.016, 291.4324, 290.215, 290.6821, 287.15, 
    287.1708, 287.268, 286.8406, 286.8147, 286.424, 286.7719, 286.9198, 
    287.2964, 287.5183, 287.7295, 288.1938, 288.709, 289.4293, 289.9579, 
    290.3052, 290.0924, 290.2802, 290.0702, 289.9719, 291.0647, 290.4507, 
    291.3725, 291.3216, 290.9042, 291.3274, 287.1855, 287.0657, 286.649, 
    286.9751, 286.3815, 286.7134, 286.904, 287.6407, 287.8032, 287.9529, 
    288.249, 288.6269, 289.2889, 289.8758, 290.4026, 290.3641, 290.3776, 
    290.4951, 290.2038, 290.5429, 290.5995, 290.451, 291.3148, 291.068, 
    291.3205, 291.1599, 287.1047, 287.3062, 287.1974, 287.4019, 287.2576, 
    287.8983, 288.0904, 288.9854, 288.6193, 289.2028, 288.6788, 288.7715, 
    289.2206, 288.7073, 289.8435, 289.0688, 290.4996, 289.7243, 290.5475, 
    290.4004, 290.6442, 290.8623, 291.1373, 291.644, 291.5267, 291.951, 
    287.6066, 287.8674, 287.845, 288.1184, 288.3198, 288.7558, 289.4538, 
    289.1916, 289.6736, 289.7702, 289.0382, 289.4871, 288.0424, 288.2762, 
    288.1376, 287.6268, 289.2513, 288.4193, 289.9664, 289.5053, 290.8311, 
    290.1764, 291.4621, 292.0106, 292.5294, 293.133, 288.0104, 287.8331, 
    288.1511, 288.5878, 288.9939, 289.5327, 289.5881, 289.6888, 289.9613, 
    290.1812, 289.7202, 290.2364, 288.3291, 289.3237, 287.7655, 288.2359, 
    288.5623, 288.4198, 289.1618, 289.3363, 290.0563, 289.6791, 291.8747, 
    290.9077, 293.5944, 292.8429, 287.771, 288.0101, 288.8374, 288.4445, 
    289.5689, 289.8561, 290.0814, 290.3686, 290.4, 290.5703, 290.2912, 
    290.5595, 289.5338, 289.998, 288.7436, 289.0461, 288.9072, 288.7543, 
    289.2259, 289.7271, 289.7387, 289.9101, 290.3614, 289.5735, 291.9979, 
    290.5053, 288.2703, 288.7267, 288.793, 288.6161, 289.8176, 289.3823, 
    290.5663, 290.2492, 290.769, 290.5106, 290.4725, 290.141, 289.9344, 
    289.402, 288.9779, 288.6418, 288.7201, 289.0892, 289.758, 290.4025, 
    290.2635, 290.7295, 289.4874, 290.0138, 289.8034, 290.335, 289.1845, 
    290.163, 288.9367, 289.0435, 289.3736, 290.0482, 290.1964, 290.3532, 
    290.2567, 289.7752, 289.6985, 289.3658, 289.2736, 289.0203, 288.8101, 
    289.0019, 289.2032, 289.7757, 290.3023, 290.8653, 291.0034, 291.6593, 
    291.1242, 292.0061, 291.2545, 292.5566, 290.2204, 291.2341, 289.3889, 
    289.5866, 289.9541, 290.7747, 290.3325, 290.85, 289.6955, 289.1015, 
    288.9488, 288.6621, 288.9554, 288.9316, 289.2121, 289.122, 289.7948, 
    289.4334, 290.4713, 290.8462, 291.9062, 292.5557, 293.2185, 293.5107, 
    293.5997, 293.6369 ;

 FSH_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSH_V =
  -13.10316, -13.10416, -13.10397, -13.10477, -13.10433, -13.10485, 
    -13.10337, -13.10419, -13.10368, -13.10326, -13.10628, -13.1048, 
    -13.10787, -13.10693, -13.1093, -13.10771, -13.10963, -13.10928, 
    -13.11039, -13.11007, -13.11147, -13.11054, -13.11223, -13.11126, 
    -13.1114, -13.11051, -13.10512, -13.1061, -13.10506, -13.1052, -13.10514, 
    -13.10434, -13.10392, -13.1031, -13.10325, -13.10386, -13.10526, 
    -13.1048, -13.10601, -13.10598, -13.10728, -13.1067, -13.10889, 
    -13.10828, -13.11009, -13.10963, -13.11006, -13.10993, -13.11007, 
    -13.10939, -13.10968, -13.10909, -13.1068, -13.10747, -13.10545, 
    -13.10419, -13.10341, -13.10283, -13.10291, -13.10307, -13.10386, 
    -13.10463, -13.10521, -13.10559, -13.10598, -13.10706, -13.10767, 
    -13.10901, -13.10878, -13.10918, -13.10958, -13.11024, -13.11013, 
    -13.11042, -13.10918, -13.11, -13.10866, -13.10901, -13.10601, -13.10493, 
    -13.10441, -13.10401, -13.10298, -13.10368, -13.1034, -13.10408, 
    -13.10451, -13.1043, -13.10561, -13.10509, -13.10771, -13.10659, 
    -13.10953, -13.10883, -13.10971, -13.10926, -13.11002, -13.10934, 
    -13.11053, -13.11078, -13.11061, -13.1113, -13.1093, -13.11006, 
    -13.10429, -13.10433, -13.10449, -13.10377, -13.10373, -13.10309, 
    -13.10367, -13.10391, -13.10454, -13.1049, -13.10525, -13.10602, 
    -13.10685, -13.10802, -13.10887, -13.10945, -13.1091, -13.10941, 
    -13.10906, -13.1089, -13.11068, -13.10968, -13.1112, -13.11112, 
    -13.11042, -13.11113, -13.10435, -13.10416, -13.10346, -13.10401, 
    -13.10302, -13.10357, -13.10387, -13.10509, -13.10538, -13.10562, 
    -13.10611, -13.10673, -13.1078, -13.10873, -13.10961, -13.10954, 
    -13.10957, -13.10976, -13.10928, -13.10983, -13.10992, -13.10968, 
    -13.11111, -13.1107, -13.11112, -13.11085, -13.10422, -13.10455, 
    -13.10437, -13.1047, -13.10446, -13.10551, -13.10583, -13.10729, 
    -13.10671, -13.10766, -13.10681, -13.10696, -13.10766, -13.10686, 
    -13.10867, -13.10742, -13.10976, -13.10848, -13.10984, -13.1096, 
    -13.11001, -13.11036, -13.11081, -13.11164, -13.11145, -13.11216, 
    -13.10505, -13.10547, -13.10545, -13.1059, -13.10622, -13.10694, 
    -13.10807, -13.10765, -13.10844, -13.10859, -13.1074, -13.10812, 
    -13.10576, -13.10614, -13.10593, -13.10507, -13.10773, -13.10637, 
    -13.10889, -13.10816, -13.11031, -13.10922, -13.11135, -13.11223, 
    -13.11312, -13.1141, -13.10572, -13.10543, -13.10596, -13.10665, 
    -13.10732, -13.1082, -13.1083, -13.10846, -13.10888, -13.10924, -13.1085, 
    -13.10933, -13.1062, -13.10785, -13.10531, -13.10607, -13.10661, 
    -13.10639, -13.10761, -13.10789, -13.10903, -13.10845, -13.112, 
    -13.11041, -13.1149, -13.11363, -13.10532, -13.10572, -13.10706, 
    -13.10643, -13.10827, -13.10871, -13.10908, -13.10954, -13.1096, 
    -13.10988, -13.10942, -13.10986, -13.1082, -13.10894, -13.10692, 
    -13.10741, -13.10719, -13.10694, -13.10771, -13.10851, -13.10854, 
    -13.10879, -13.10947, -13.10827, -13.11217, -13.10971, -13.10615, 
    -13.10687, -13.107, -13.10671, -13.10867, -13.10796, -13.10987, 
    -13.10935, -13.11021, -13.10978, -13.10972, -13.10918, -13.10884, 
    -13.10799, -13.1073, -13.10676, -13.10688, -13.10748, -13.10856, 
    -13.1096, -13.10937, -13.11014, -13.10813, -13.10896, -13.10864, 
    -13.10949, -13.10763, -13.10915, -13.10724, -13.10741, -13.10794, 
    -13.109, -13.10927, -13.10952, -13.10937, -13.10859, -13.10847, 
    -13.10793, -13.10778, -13.10737, -13.10703, -13.10734, -13.10766, 
    -13.1086, -13.10943, -13.11036, -13.11059, -13.11164, -13.11076, 
    -13.11218, -13.11093, -13.11312, -13.10927, -13.11093, -13.10797, 
    -13.1083, -13.10885, -13.11019, -13.10949, -13.11032, -13.10847, 
    -13.10749, -13.10726, -13.10679, -13.10727, -13.10723, -13.10769, 
    -13.10754, -13.10863, -13.10805, -13.10971, -13.11032, -13.11207, 
    -13.11315, -13.11427, -13.11476, -13.11491, -13.11498 ;

 FSM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSNO_EFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSR =
  1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 1.049531, 
    1.049531, 1.049531 ;

 FSRND =
  0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 0.1566151, 
    0.1566151, 0.1566151 ;

 FSRNDLN =
  0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372 ;

 FSRNI =
  0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 0.3681505, 
    0.3681505, 0.3681505 ;

 FSRVD =
  0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 0.09373803, 
    0.09373803, 0.09373803 ;

 FSRVDLN =
  0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678 ;

 FSRVI =
  0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 0.4310275, 
    0.4310275, 0.4310275 ;

 FUELC =
  0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806 ;

 F_DENIT =
  2.809608e-14, 2.822132e-14, 2.81969e-14, 2.8298e-14, 2.824186e-14, 
    2.830805e-14, 2.812131e-14, 2.822615e-14, 2.815916e-14, 2.81071e-14, 
    2.849427e-14, 2.830232e-14, 2.869362e-14, 2.857102e-14, 2.887894e-14, 
    2.867451e-14, 2.892015e-14, 2.887291e-14, 2.901485e-14, 2.897413e-14, 
    2.91559e-14, 2.903356e-14, 2.925006e-14, 2.91266e-14, 2.91459e-14, 
    2.902941e-14, 2.834104e-14, 2.847056e-14, 2.833334e-14, 2.83518e-14, 
    2.834347e-14, 2.824293e-14, 2.819234e-14, 2.808624e-14, 2.810545e-14, 
    2.818333e-14, 2.835992e-14, 2.829987e-14, 2.845101e-14, 2.84476e-14, 
    2.861606e-14, 2.854006e-14, 2.882346e-14, 2.874281e-14, 2.89758e-14, 
    2.891714e-14, 2.897301e-14, 2.895601e-14, 2.897315e-14, 2.88872e-14, 
    2.892397e-14, 2.884833e-14, 2.85546e-14, 2.864101e-14, 2.838332e-14, 
    2.822863e-14, 2.812581e-14, 2.805297e-14, 2.806321e-14, 2.808286e-14, 
    2.818374e-14, 2.827859e-14, 2.835094e-14, 2.839934e-14, 2.844704e-14, 
    2.859176e-14, 2.866824e-14, 2.883974e-14, 2.880871e-14, 2.886118e-14, 
    2.891128e-14, 2.899547e-14, 2.898159e-14, 2.901868e-14, 2.885963e-14, 
    2.896532e-14, 2.879083e-14, 2.883854e-14, 2.846047e-14, 2.831616e-14, 
    2.825504e-14, 2.820137e-14, 2.807112e-14, 2.816105e-14, 2.812557e-14, 
    2.820984e-14, 2.826346e-14, 2.823689e-14, 2.840064e-14, 2.833692e-14, 
    2.867274e-14, 2.8528e-14, 2.890547e-14, 2.881501e-14, 2.892707e-14, 
    2.886986e-14, 2.896786e-14, 2.887962e-14, 2.903243e-14, 2.906577e-14, 
    2.904294e-14, 2.913036e-14, 2.887457e-14, 2.897278e-14, 2.82363e-14, 
    2.824063e-14, 2.826075e-14, 2.817219e-14, 2.816675e-14, 2.808558e-14, 
    2.815772e-14, 2.818848e-14, 2.826649e-14, 2.831267e-14, 2.835656e-14, 
    2.84532e-14, 2.856119e-14, 2.871226e-14, 2.882085e-14, 2.889366e-14, 
    2.884896e-14, 2.888837e-14, 2.884427e-14, 2.882356e-14, 2.905322e-14, 
    2.892423e-14, 2.911771e-14, 2.9107e-14, 2.901938e-14, 2.910813e-14, 
    2.824362e-14, 2.821868e-14, 2.813231e-14, 2.819985e-14, 2.807669e-14, 
    2.814563e-14, 2.818527e-14, 2.833826e-14, 2.837182e-14, 2.840305e-14, 
    2.846465e-14, 2.854377e-14, 2.868271e-14, 2.880364e-14, 2.891409e-14, 
    2.890595e-14, 2.890879e-14, 2.893346e-14, 2.887228e-14, 2.894345e-14, 
    2.895539e-14, 2.892413e-14, 2.910549e-14, 2.905365e-14, 2.910667e-14, 
    2.907286e-14, 2.822674e-14, 2.82686e-14, 2.824593e-14, 2.828852e-14, 
    2.825848e-14, 2.839191e-14, 2.84319e-14, 2.861922e-14, 2.854222e-14, 
    2.866468e-14, 2.855459e-14, 2.85741e-14, 2.866868e-14, 2.856045e-14, 
    2.879692e-14, 2.86366e-14, 2.893439e-14, 2.877425e-14, 2.894438e-14, 
    2.891341e-14, 2.896458e-14, 2.901049e-14, 2.906815e-14, 2.917476e-14, 
    2.915e-14, 2.923916e-14, 2.833103e-14, 2.838539e-14, 2.838055e-14, 
    2.843742e-14, 2.847951e-14, 2.857078e-14, 2.871728e-14, 2.866211e-14, 
    2.876326e-14, 2.87836e-14, 2.862981e-14, 2.872423e-14, 2.842152e-14, 
    2.847038e-14, 2.844123e-14, 2.833496e-14, 2.867466e-14, 2.850022e-14, 
    2.882235e-14, 2.872773e-14, 2.900387e-14, 2.886652e-14, 2.91364e-14, 
    2.925202e-14, 2.936066e-14, 2.948791e-14, 2.841501e-14, 2.837801e-14, 
    2.844413e-14, 2.853579e-14, 2.86207e-14, 2.87338e-14, 2.874532e-14, 
    2.876649e-14, 2.882135e-14, 2.886755e-14, 2.877317e-14, 2.887905e-14, 
    2.848178e-14, 2.868978e-14, 2.836375e-14, 2.84619e-14, 2.853002e-14, 
    2.850008e-14, 2.865548e-14, 2.869211e-14, 2.884117e-14, 2.876407e-14, 
    2.922344e-14, 2.902005e-14, 2.95847e-14, 2.942677e-14, 2.836508e-14, 
    2.841476e-14, 2.858796e-14, 2.850551e-14, 2.874126e-14, 2.879937e-14, 
    2.884654e-14, 2.890698e-14, 2.891343e-14, 2.894924e-14, 2.889051e-14, 
    2.894686e-14, 2.873377e-14, 2.882894e-14, 2.856783e-14, 2.863132e-14, 
    2.860207e-14, 2.856999e-14, 2.866887e-14, 2.877439e-14, 2.877655e-14, 
    2.881037e-14, 2.890591e-14, 2.874176e-14, 2.924972e-14, 2.893592e-14, 
    2.846897e-14, 2.856487e-14, 2.857847e-14, 2.854132e-14, 2.879348e-14, 
    2.870206e-14, 2.894836e-14, 2.88817e-14, 2.899082e-14, 2.893659e-14, 
    2.892856e-14, 2.885891e-14, 2.881552e-14, 2.870607e-14, 2.861699e-14, 
    2.854641e-14, 2.856276e-14, 2.864032e-14, 2.878076e-14, 2.891373e-14, 
    2.888458e-14, 2.898221e-14, 2.872365e-14, 2.883205e-14, 2.879011e-14, 
    2.889933e-14, 2.866056e-14, 2.886451e-14, 2.860846e-14, 2.863084e-14, 
    2.870018e-14, 2.883982e-14, 2.887058e-14, 2.890361e-14, 2.888316e-14, 
    2.87845e-14, 2.876828e-14, 2.869831e-14, 2.867901e-14, 2.862573e-14, 
    2.858161e-14, 2.862189e-14, 2.866416e-14, 2.878432e-14, 2.889267e-14, 
    2.901084e-14, 2.903975e-14, 2.91781e-14, 2.906551e-14, 2.925136e-14, 
    2.909343e-14, 2.936677e-14, 2.887617e-14, 2.908917e-14, 2.870332e-14, 
    2.874479e-14, 2.881995e-14, 2.899231e-14, 2.889912e-14, 2.900805e-14, 
    2.876762e-14, 2.864306e-14, 2.861075e-14, 2.855067e-14, 2.861208e-14, 
    2.860708e-14, 2.866588e-14, 2.864693e-14, 2.878824e-14, 2.87123e-14, 
    2.892804e-14, 2.900687e-14, 2.922955e-14, 2.936619e-14, 2.95053e-14, 
    2.956674e-14, 2.958544e-14, 2.959324e-14 ;

 F_DENIT_vr =
  1.604315e-12, 1.611466e-12, 1.610072e-12, 1.615845e-12, 1.612639e-12, 
    1.616419e-12, 1.605756e-12, 1.611742e-12, 1.607917e-12, 1.604944e-12, 
    1.627052e-12, 1.616091e-12, 1.638435e-12, 1.631435e-12, 1.649017e-12, 
    1.637344e-12, 1.65137e-12, 1.648673e-12, 1.656778e-12, 1.654453e-12, 
    1.664832e-12, 1.657846e-12, 1.670208e-12, 1.663159e-12, 1.664261e-12, 
    1.657609e-12, 1.618303e-12, 1.625698e-12, 1.617863e-12, 1.618917e-12, 
    1.618441e-12, 1.612701e-12, 1.609812e-12, 1.603753e-12, 1.60485e-12, 
    1.609297e-12, 1.619381e-12, 1.615952e-12, 1.624582e-12, 1.624387e-12, 
    1.634006e-12, 1.629667e-12, 1.645849e-12, 1.641244e-12, 1.654548e-12, 
    1.651199e-12, 1.654389e-12, 1.653418e-12, 1.654397e-12, 1.649489e-12, 
    1.651589e-12, 1.64727e-12, 1.630497e-12, 1.635431e-12, 1.620717e-12, 
    1.611884e-12, 1.606013e-12, 1.601854e-12, 1.602438e-12, 1.60356e-12, 
    1.609321e-12, 1.614737e-12, 1.618868e-12, 1.621632e-12, 1.624355e-12, 
    1.632619e-12, 1.636986e-12, 1.646779e-12, 1.645007e-12, 1.648003e-12, 
    1.650864e-12, 1.655671e-12, 1.654879e-12, 1.656997e-12, 1.647915e-12, 
    1.65395e-12, 1.643986e-12, 1.64671e-12, 1.625122e-12, 1.616882e-12, 
    1.613392e-12, 1.610328e-12, 1.60289e-12, 1.608025e-12, 1.605999e-12, 
    1.610811e-12, 1.613873e-12, 1.612356e-12, 1.621706e-12, 1.618068e-12, 
    1.637243e-12, 1.628978e-12, 1.650532e-12, 1.645367e-12, 1.651765e-12, 
    1.648499e-12, 1.654095e-12, 1.649056e-12, 1.657782e-12, 1.659685e-12, 
    1.658382e-12, 1.663374e-12, 1.648768e-12, 1.654375e-12, 1.612322e-12, 
    1.612569e-12, 1.613718e-12, 1.608661e-12, 1.60835e-12, 1.603715e-12, 
    1.607835e-12, 1.609592e-12, 1.614046e-12, 1.616682e-12, 1.619189e-12, 
    1.624707e-12, 1.630873e-12, 1.639499e-12, 1.6457e-12, 1.649858e-12, 
    1.647305e-12, 1.649556e-12, 1.647038e-12, 1.645855e-12, 1.658969e-12, 
    1.651604e-12, 1.662652e-12, 1.66204e-12, 1.657036e-12, 1.662104e-12, 
    1.61274e-12, 1.611316e-12, 1.606384e-12, 1.610241e-12, 1.603208e-12, 
    1.607145e-12, 1.609408e-12, 1.618144e-12, 1.620061e-12, 1.621844e-12, 
    1.625361e-12, 1.629879e-12, 1.637812e-12, 1.644717e-12, 1.651024e-12, 
    1.65056e-12, 1.650722e-12, 1.65213e-12, 1.648637e-12, 1.652701e-12, 
    1.653383e-12, 1.651597e-12, 1.661954e-12, 1.658993e-12, 1.662021e-12, 
    1.660091e-12, 1.611776e-12, 1.614166e-12, 1.612872e-12, 1.615303e-12, 
    1.613588e-12, 1.621207e-12, 1.623491e-12, 1.634187e-12, 1.62979e-12, 
    1.636783e-12, 1.630496e-12, 1.631611e-12, 1.637011e-12, 1.630831e-12, 
    1.644334e-12, 1.63518e-12, 1.652184e-12, 1.64304e-12, 1.652754e-12, 
    1.650985e-12, 1.653907e-12, 1.656529e-12, 1.659821e-12, 1.665909e-12, 
    1.664495e-12, 1.669586e-12, 1.617731e-12, 1.620835e-12, 1.620559e-12, 
    1.623806e-12, 1.626209e-12, 1.631421e-12, 1.639786e-12, 1.636636e-12, 
    1.642412e-12, 1.643573e-12, 1.634792e-12, 1.640183e-12, 1.622898e-12, 
    1.625688e-12, 1.624023e-12, 1.617956e-12, 1.637353e-12, 1.627392e-12, 
    1.645786e-12, 1.640383e-12, 1.656151e-12, 1.648308e-12, 1.663718e-12, 
    1.67032e-12, 1.676524e-12, 1.68379e-12, 1.622527e-12, 1.620414e-12, 
    1.624189e-12, 1.629423e-12, 1.634272e-12, 1.64073e-12, 1.641388e-12, 
    1.642596e-12, 1.645729e-12, 1.648367e-12, 1.642978e-12, 1.649024e-12, 
    1.626339e-12, 1.638216e-12, 1.619599e-12, 1.625204e-12, 1.629094e-12, 
    1.627384e-12, 1.636258e-12, 1.638349e-12, 1.646861e-12, 1.642458e-12, 
    1.668688e-12, 1.657075e-12, 1.689317e-12, 1.680299e-12, 1.619675e-12, 
    1.622512e-12, 1.632402e-12, 1.627694e-12, 1.641156e-12, 1.644474e-12, 
    1.647167e-12, 1.650619e-12, 1.650986e-12, 1.653032e-12, 1.649678e-12, 
    1.652896e-12, 1.640728e-12, 1.646162e-12, 1.631253e-12, 1.634878e-12, 
    1.633208e-12, 1.631376e-12, 1.637022e-12, 1.643047e-12, 1.643171e-12, 
    1.645102e-12, 1.650557e-12, 1.641184e-12, 1.670189e-12, 1.652271e-12, 
    1.625608e-12, 1.631084e-12, 1.63186e-12, 1.629739e-12, 1.644137e-12, 
    1.638917e-12, 1.652981e-12, 1.649175e-12, 1.655406e-12, 1.652309e-12, 
    1.65185e-12, 1.647873e-12, 1.645396e-12, 1.639146e-12, 1.63406e-12, 
    1.630029e-12, 1.630963e-12, 1.635392e-12, 1.643411e-12, 1.651004e-12, 
    1.649339e-12, 1.654914e-12, 1.64015e-12, 1.64634e-12, 1.643945e-12, 
    1.650182e-12, 1.636548e-12, 1.648193e-12, 1.633573e-12, 1.634851e-12, 
    1.63881e-12, 1.646784e-12, 1.64854e-12, 1.650426e-12, 1.649258e-12, 
    1.643625e-12, 1.642698e-12, 1.638703e-12, 1.637601e-12, 1.634559e-12, 
    1.632039e-12, 1.63434e-12, 1.636753e-12, 1.643614e-12, 1.649801e-12, 
    1.656549e-12, 1.658199e-12, 1.666099e-12, 1.659671e-12, 1.670283e-12, 
    1.661265e-12, 1.676873e-12, 1.648859e-12, 1.661022e-12, 1.638989e-12, 
    1.641357e-12, 1.645649e-12, 1.655491e-12, 1.65017e-12, 1.65639e-12, 
    1.642661e-12, 1.635549e-12, 1.633703e-12, 1.630273e-12, 1.633779e-12, 
    1.633494e-12, 1.636851e-12, 1.635769e-12, 1.643838e-12, 1.639502e-12, 
    1.651821e-12, 1.656323e-12, 1.669037e-12, 1.67684e-12, 1.684783e-12, 
    1.688291e-12, 1.689359e-12, 1.689804e-12,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_N2O_DENIT =
  7.628954e-16, 7.636266e-16, 7.634834e-16, 7.640685e-16, 7.637434e-16, 
    7.641247e-16, 7.630404e-16, 7.636513e-16, 7.632608e-16, 7.629551e-16, 
    7.651825e-16, 7.64089e-16, 7.662893e-16, 7.656084e-16, 7.673018e-16, 
    7.661831e-16, 7.675239e-16, 7.672667e-16, 7.680303e-16, 7.678115e-16, 
    7.687777e-16, 7.681287e-16, 7.69268e-16, 7.686216e-16, 7.68723e-16, 
    7.681041e-16, 7.643143e-16, 7.650529e-16, 7.642691e-16, 7.643752e-16, 
    7.643266e-16, 7.637477e-16, 7.634549e-16, 7.62832e-16, 7.629443e-16, 
    7.634005e-16, 7.64418e-16, 7.640724e-16, 7.649331e-16, 7.649138e-16, 
    7.658568e-16, 7.654332e-16, 7.66997e-16, 7.665537e-16, 7.678199e-16, 
    7.675035e-16, 7.67804e-16, 7.677119e-16, 7.678033e-16, 7.673402e-16, 
    7.675378e-16, 7.671279e-16, 7.655209e-16, 7.660009e-16, 7.645539e-16, 
    7.63666e-16, 7.630648e-16, 7.626361e-16, 7.626955e-16, 7.628117e-16, 
    7.634018e-16, 7.639497e-16, 7.643644e-16, 7.646396e-16, 7.649092e-16, 
    7.657233e-16, 7.661455e-16, 7.670851e-16, 7.669148e-16, 7.672006e-16, 
    7.674713e-16, 7.679234e-16, 7.678486e-16, 7.680465e-16, 7.671888e-16, 
    7.677604e-16, 7.668121e-16, 7.670731e-16, 7.649937e-16, 7.641684e-16, 
    7.638179e-16, 7.635051e-16, 7.627418e-16, 7.632698e-16, 7.630615e-16, 
    7.635517e-16, 7.638619e-16, 7.637073e-16, 7.646463e-16, 7.642822e-16, 
    7.661695e-16, 7.653644e-16, 7.674406e-16, 7.669482e-16, 7.675556e-16, 
    7.67246e-16, 7.677745e-16, 7.67298e-16, 7.681186e-16, 7.682965e-16, 
    7.681737e-16, 7.686366e-16, 7.672674e-16, 7.677979e-16, 7.637071e-16, 
    7.637324e-16, 7.638478e-16, 7.63334e-16, 7.633019e-16, 7.628252e-16, 
    7.632473e-16, 7.63427e-16, 7.638777e-16, 7.641429e-16, 7.643936e-16, 
    7.649427e-16, 7.655491e-16, 7.663847e-16, 7.669794e-16, 7.673742e-16, 
    7.671313e-16, 7.673446e-16, 7.671049e-16, 7.66991e-16, 7.682283e-16, 
    7.675374e-16, 7.685684e-16, 7.685118e-16, 7.680462e-16, 7.685163e-16, 
    7.637486e-16, 7.636032e-16, 7.631e-16, 7.634929e-16, 7.627717e-16, 
    7.631767e-16, 7.634077e-16, 7.642898e-16, 7.644801e-16, 7.646582e-16, 
    7.650061e-16, 7.654499e-16, 7.662215e-16, 7.668845e-16, 7.674841e-16, 
    7.674393e-16, 7.674545e-16, 7.67587e-16, 7.672558e-16, 7.676398e-16, 
    7.677037e-16, 7.67535e-16, 7.685023e-16, 7.682276e-16, 7.68508e-16, 
    7.683281e-16, 7.636493e-16, 7.638906e-16, 7.63759e-16, 7.64005e-16, 
    7.638308e-16, 7.645963e-16, 7.648228e-16, 7.658719e-16, 7.654414e-16, 
    7.661226e-16, 7.655093e-16, 7.656186e-16, 7.661443e-16, 7.655405e-16, 
    7.668468e-16, 7.659645e-16, 7.675914e-16, 7.667215e-16, 7.676442e-16, 
    7.674761e-16, 7.67751e-16, 7.679974e-16, 7.683031e-16, 7.688663e-16, 
    7.687349e-16, 7.692013e-16, 7.642488e-16, 7.645589e-16, 7.645305e-16, 
    7.648528e-16, 7.650899e-16, 7.656014e-16, 7.664116e-16, 7.661068e-16, 
    7.666622e-16, 7.667741e-16, 7.659262e-16, 7.664476e-16, 7.647587e-16, 
    7.650349e-16, 7.648691e-16, 7.642636e-16, 7.661726e-16, 7.652007e-16, 
    7.669815e-16, 7.664616e-16, 7.679606e-16, 7.672212e-16, 7.686629e-16, 
    7.692693e-16, 7.69828e-16, 7.704768e-16, 7.647263e-16, 7.645148e-16, 
    7.648895e-16, 7.654065e-16, 7.658778e-16, 7.665014e-16, 7.665637e-16, 
    7.666795e-16, 7.669789e-16, 7.672306e-16, 7.667156e-16, 7.672915e-16, 
    7.650999e-16, 7.662554e-16, 7.64427e-16, 7.649852e-16, 7.653665e-16, 
    7.651982e-16, 7.660631e-16, 7.662644e-16, 7.670815e-16, 7.666591e-16, 
    7.691192e-16, 7.680456e-16, 7.709612e-16, 7.701652e-16, 7.644405e-16, 
    7.647224e-16, 7.656959e-16, 7.652345e-16, 7.665405e-16, 7.668599e-16, 
    7.671158e-16, 7.674444e-16, 7.674777e-16, 7.676711e-16, 7.673526e-16, 
    7.67657e-16, 7.664956e-16, 7.670172e-16, 7.655771e-16, 7.659298e-16, 
    7.657667e-16, 7.655873e-16, 7.661353e-16, 7.667165e-16, 7.667267e-16, 
    7.669115e-16, 7.67434e-16, 7.665335e-16, 7.692561e-16, 7.675936e-16, 
    7.650285e-16, 7.655671e-16, 7.656411e-16, 7.654335e-16, 7.668261e-16, 
    7.663244e-16, 7.676662e-16, 7.673052e-16, 7.678925e-16, 7.676014e-16, 
    7.67557e-16, 7.671798e-16, 7.669424e-16, 7.663424e-16, 7.658493e-16, 
    7.654556e-16, 7.655459e-16, 7.659777e-16, 7.667497e-16, 7.674732e-16, 
    7.67315e-16, 7.678397e-16, 7.664332e-16, 7.670279e-16, 7.667977e-16, 
    7.673919e-16, 7.660962e-16, 7.672173e-16, 7.658067e-16, 7.659301e-16, 
    7.663125e-16, 7.67079e-16, 7.672438e-16, 7.674233e-16, 7.673109e-16, 
    7.66774e-16, 7.666839e-16, 7.662985e-16, 7.661919e-16, 7.65897e-16, 
    7.656506e-16, 7.658749e-16, 7.661081e-16, 7.667684e-16, 7.673583e-16, 
    7.67993e-16, 7.681465e-16, 7.68879e-16, 7.682843e-16, 7.692621e-16, 
    7.684338e-16, 7.698557e-16, 7.672778e-16, 7.684199e-16, 7.663295e-16, 
    7.665563e-16, 7.669693e-16, 7.679007e-16, 7.673972e-16, 7.679841e-16, 
    7.666799e-16, 7.659943e-16, 7.658134e-16, 7.65479e-16, 7.658197e-16, 
    7.657921e-16, 7.661169e-16, 7.660114e-16, 7.667883e-16, 7.663713e-16, 
    7.675474e-16, 7.679713e-16, 7.691456e-16, 7.698516e-16, 7.705578e-16, 
    7.708659e-16, 7.709592e-16, 7.709976e-16 ;

 F_N2O_NIT =
  2.408731e-14, 2.429515e-14, 2.425467e-14, 2.442284e-14, 2.432947e-14, 
    2.44397e-14, 2.412936e-14, 2.430341e-14, 2.419222e-14, 2.410595e-14, 
    2.475091e-14, 2.443034e-14, 2.508615e-14, 2.488003e-14, 2.539948e-14, 
    2.505402e-14, 2.546943e-14, 2.538947e-14, 2.56305e-14, 2.556132e-14, 
    2.587092e-14, 2.566245e-14, 2.603216e-14, 2.582105e-14, 2.585402e-14, 
    2.565558e-14, 2.449469e-14, 2.47109e-14, 2.448191e-14, 2.451267e-14, 
    2.449886e-14, 2.433139e-14, 2.424723e-14, 2.407143e-14, 2.410329e-14, 
    2.423243e-14, 2.452649e-14, 2.442646e-14, 2.467895e-14, 2.467323e-14, 
    2.495588e-14, 2.482823e-14, 2.530578e-14, 2.516957e-14, 2.556421e-14, 
    2.546466e-14, 2.555952e-14, 2.553073e-14, 2.555989e-14, 2.541398e-14, 
    2.547644e-14, 2.534823e-14, 2.485214e-14, 2.499743e-14, 2.45654e-14, 
    2.43075e-14, 2.413697e-14, 2.401634e-14, 2.403337e-14, 2.406586e-14, 
    2.423318e-14, 2.439104e-14, 2.45117e-14, 2.459258e-14, 2.46724e-14, 
    2.491487e-14, 2.504369e-14, 2.533337e-14, 2.528095e-14, 2.536977e-14, 
    2.545476e-14, 2.559779e-14, 2.557422e-14, 2.563734e-14, 2.536741e-14, 
    2.554664e-14, 2.525111e-14, 2.533176e-14, 2.469418e-14, 2.445343e-14, 
    2.435149e-14, 2.426243e-14, 2.404647e-14, 2.41955e-14, 2.413669e-14, 
    2.42767e-14, 2.436589e-14, 2.432175e-14, 2.459479e-14, 2.448845e-14, 
    2.505133e-14, 2.480807e-14, 2.544484e-14, 2.52917e-14, 2.548161e-14, 
    2.538461e-14, 2.555093e-14, 2.540122e-14, 2.566084e-14, 2.571756e-14, 
    2.567879e-14, 2.582786e-14, 2.539291e-14, 2.55595e-14, 2.432053e-14, 
    2.432773e-14, 2.436126e-14, 2.421403e-14, 2.420504e-14, 2.407054e-14, 
    2.419019e-14, 2.424124e-14, 2.437106e-14, 2.444802e-14, 2.452129e-14, 
    2.468281e-14, 2.486383e-14, 2.511811e-14, 2.530161e-14, 2.5425e-14, 
    2.53493e-14, 2.541612e-14, 2.534142e-14, 2.530644e-14, 2.569629e-14, 
    2.547701e-14, 2.580639e-14, 2.57881e-14, 2.563882e-14, 2.579015e-14, 
    2.433278e-14, 2.429138e-14, 2.414795e-14, 2.426016e-14, 2.405592e-14, 
    2.417013e-14, 2.423593e-14, 2.449067e-14, 2.454682e-14, 2.459895e-14, 
    2.470207e-14, 2.483474e-14, 2.506837e-14, 2.527255e-14, 2.54597e-14, 
    2.544596e-14, 2.545079e-14, 2.549269e-14, 2.538897e-14, 2.550973e-14, 
    2.553003e-14, 2.547697e-14, 2.578565e-14, 2.569726e-14, 2.57877e-14, 
    2.573013e-14, 2.430483e-14, 2.437451e-14, 2.433684e-14, 2.44077e-14, 
    2.435777e-14, 2.458021e-14, 2.46471e-14, 2.496135e-14, 2.483212e-14, 
    2.503795e-14, 2.485298e-14, 2.488571e-14, 2.504468e-14, 2.486295e-14, 
    2.526127e-14, 2.499087e-14, 2.549432e-14, 2.522301e-14, 2.551136e-14, 
    2.545887e-14, 2.55458e-14, 2.562379e-14, 2.572208e-14, 2.590396e-14, 
    2.586178e-14, 2.601426e-14, 2.447859e-14, 2.456934e-14, 2.456133e-14, 
    2.465646e-14, 2.472694e-14, 2.488005e-14, 2.512664e-14, 2.503376e-14, 
    2.52044e-14, 2.523873e-14, 2.497953e-14, 2.513851e-14, 2.463014e-14, 
    2.471191e-14, 2.46632e-14, 2.448571e-14, 2.505513e-14, 2.476206e-14, 
    2.530462e-14, 2.514481e-14, 2.561266e-14, 2.537943e-14, 2.583857e-14, 
    2.603616e-14, 2.622282e-14, 2.644184e-14, 2.461893e-14, 2.455718e-14, 
    2.466778e-14, 2.482124e-14, 2.496405e-14, 2.515458e-14, 2.517411e-14, 
    2.520989e-14, 2.530272e-14, 2.538091e-14, 2.522121e-14, 2.540052e-14, 
    2.47309e-14, 2.508065e-14, 2.453383e-14, 2.469784e-14, 2.481214e-14, 
    2.476196e-14, 2.502312e-14, 2.508488e-14, 2.533666e-14, 2.520634e-14, 
    2.598732e-14, 2.564027e-14, 2.660922e-14, 2.633657e-14, 2.453563e-14, 
    2.46187e-14, 2.490898e-14, 2.477065e-14, 2.516731e-14, 2.526545e-14, 
    2.534537e-14, 2.544773e-14, 2.545879e-14, 2.551955e-14, 2.542001e-14, 
    2.551561e-14, 2.515496e-14, 2.531579e-14, 2.487568e-14, 2.498243e-14, 
    2.493329e-14, 2.487944e-14, 2.504581e-14, 2.52237e-14, 2.52275e-14, 
    2.528467e-14, 2.544618e-14, 2.516888e-14, 2.603229e-14, 2.54973e-14, 
    2.470946e-14, 2.487021e-14, 2.48932e-14, 2.483084e-14, 2.52556e-14, 
    2.510126e-14, 2.551807e-14, 2.540506e-14, 2.559035e-14, 2.549819e-14, 
    2.548464e-14, 2.536656e-14, 2.529318e-14, 2.510831e-14, 2.495839e-14, 
    2.483984e-14, 2.486738e-14, 2.499769e-14, 2.523459e-14, 2.545976e-14, 
    2.541035e-14, 2.557621e-14, 2.513839e-14, 2.53215e-14, 2.525065e-14, 
    2.54356e-14, 2.503129e-14, 2.537544e-14, 2.494371e-14, 2.49814e-14, 
    2.509819e-14, 2.533399e-14, 2.538629e-14, 2.544222e-14, 2.54077e-14, 
    2.524064e-14, 2.521331e-14, 2.509533e-14, 2.506281e-14, 2.497317e-14, 
    2.489907e-14, 2.496676e-14, 2.503795e-14, 2.524068e-14, 2.542411e-14, 
    2.562487e-14, 2.567413e-14, 2.590999e-14, 2.571791e-14, 2.603528e-14, 
    2.576534e-14, 2.623353e-14, 2.539544e-14, 2.575746e-14, 2.510351e-14, 
    2.517354e-14, 2.530047e-14, 2.559282e-14, 2.543476e-14, 2.561965e-14, 
    2.521224e-14, 2.50022e-14, 2.4948e-14, 2.484704e-14, 2.49503e-14, 
    2.494189e-14, 2.504089e-14, 2.500905e-14, 2.524742e-14, 2.511923e-14, 
    2.548427e-14, 2.561816e-14, 2.599823e-14, 2.623265e-14, 2.64724e-14, 
    2.65786e-14, 2.661096e-14, 2.66245e-14 ;

 F_NIT =
  4.014551e-11, 4.049193e-11, 4.042445e-11, 4.070474e-11, 4.054912e-11, 
    4.073283e-11, 4.021559e-11, 4.050569e-11, 4.032037e-11, 4.017659e-11, 
    4.125151e-11, 4.071723e-11, 4.181026e-11, 4.146671e-11, 4.233246e-11, 
    4.17567e-11, 4.244905e-11, 4.231578e-11, 4.27175e-11, 4.260221e-11, 
    4.31182e-11, 4.277076e-11, 4.338693e-11, 4.303508e-11, 4.309002e-11, 
    4.27593e-11, 4.082448e-11, 4.118484e-11, 4.080318e-11, 4.085445e-11, 
    4.083144e-11, 4.055232e-11, 4.041205e-11, 4.011905e-11, 4.017215e-11, 
    4.038738e-11, 4.087749e-11, 4.071076e-11, 4.113158e-11, 4.112206e-11, 
    4.159313e-11, 4.138039e-11, 4.21763e-11, 4.194928e-11, 4.260701e-11, 
    4.24411e-11, 4.25992e-11, 4.255122e-11, 4.259982e-11, 4.235663e-11, 
    4.246073e-11, 4.224705e-11, 4.142024e-11, 4.166238e-11, 4.094233e-11, 
    4.05125e-11, 4.022828e-11, 4.002723e-11, 4.005561e-11, 4.010977e-11, 
    4.038864e-11, 4.065173e-11, 4.085283e-11, 4.098763e-11, 4.112067e-11, 
    4.152479e-11, 4.173948e-11, 4.222228e-11, 4.213492e-11, 4.228295e-11, 
    4.24246e-11, 4.266299e-11, 4.26237e-11, 4.272889e-11, 4.227901e-11, 
    4.257773e-11, 4.208518e-11, 4.22196e-11, 4.115696e-11, 4.075572e-11, 
    4.058582e-11, 4.043738e-11, 4.007744e-11, 4.032583e-11, 4.022781e-11, 
    4.046117e-11, 4.060982e-11, 4.053626e-11, 4.099131e-11, 4.081408e-11, 
    4.175221e-11, 4.134678e-11, 4.240807e-11, 4.215283e-11, 4.246935e-11, 
    4.230769e-11, 4.258488e-11, 4.233536e-11, 4.276807e-11, 4.28626e-11, 
    4.279798e-11, 4.304643e-11, 4.232152e-11, 4.259916e-11, 4.053422e-11, 
    4.054622e-11, 4.06021e-11, 4.035672e-11, 4.034173e-11, 4.011757e-11, 
    4.031699e-11, 4.040206e-11, 4.061843e-11, 4.07467e-11, 4.086882e-11, 
    4.113801e-11, 4.143972e-11, 4.186352e-11, 4.216935e-11, 4.2375e-11, 
    4.224883e-11, 4.236021e-11, 4.22357e-11, 4.217741e-11, 4.282716e-11, 
    4.246168e-11, 4.301064e-11, 4.298017e-11, 4.273137e-11, 4.298359e-11, 
    4.055463e-11, 4.048563e-11, 4.024659e-11, 4.043359e-11, 4.009319e-11, 
    4.028355e-11, 4.039321e-11, 4.081778e-11, 4.091136e-11, 4.099825e-11, 
    4.117012e-11, 4.139123e-11, 4.178061e-11, 4.212092e-11, 4.243283e-11, 
    4.240993e-11, 4.241799e-11, 4.248782e-11, 4.231495e-11, 4.251622e-11, 
    4.255005e-11, 4.246162e-11, 4.297608e-11, 4.282877e-11, 4.297951e-11, 
    4.288355e-11, 4.050804e-11, 4.062419e-11, 4.05614e-11, 4.06795e-11, 
    4.059628e-11, 4.096701e-11, 4.10785e-11, 4.160226e-11, 4.138687e-11, 
    4.172991e-11, 4.142164e-11, 4.147618e-11, 4.174113e-11, 4.143826e-11, 
    4.210211e-11, 4.165145e-11, 4.249053e-11, 4.203836e-11, 4.251894e-11, 
    4.243145e-11, 4.257633e-11, 4.270632e-11, 4.287013e-11, 4.317326e-11, 
    4.310296e-11, 4.33571e-11, 4.079765e-11, 4.094889e-11, 4.093556e-11, 
    4.109411e-11, 4.121157e-11, 4.146675e-11, 4.187774e-11, 4.172293e-11, 
    4.200734e-11, 4.206455e-11, 4.163255e-11, 4.189752e-11, 4.105023e-11, 
    4.118651e-11, 4.110533e-11, 4.080952e-11, 4.175855e-11, 4.127009e-11, 
    4.217436e-11, 4.190802e-11, 4.268777e-11, 4.229906e-11, 4.306429e-11, 
    4.339361e-11, 4.370469e-11, 4.406973e-11, 4.103155e-11, 4.092864e-11, 
    4.111297e-11, 4.136873e-11, 4.160675e-11, 4.192429e-11, 4.195684e-11, 
    4.201649e-11, 4.217119e-11, 4.230151e-11, 4.203536e-11, 4.23342e-11, 
    4.121816e-11, 4.180109e-11, 4.088972e-11, 4.116307e-11, 4.135358e-11, 
    4.126994e-11, 4.170521e-11, 4.180813e-11, 4.222776e-11, 4.201057e-11, 
    4.33122e-11, 4.273379e-11, 4.434871e-11, 4.389429e-11, 4.089271e-11, 
    4.103117e-11, 4.151497e-11, 4.128441e-11, 4.194552e-11, 4.210909e-11, 
    4.224228e-11, 4.241289e-11, 4.243132e-11, 4.253259e-11, 4.236669e-11, 
    4.252602e-11, 4.192493e-11, 4.219299e-11, 4.145947e-11, 4.163739e-11, 
    4.155548e-11, 4.146574e-11, 4.174302e-11, 4.20395e-11, 4.204583e-11, 
    4.214112e-11, 4.24103e-11, 4.194813e-11, 4.338716e-11, 4.24955e-11, 
    4.118243e-11, 4.145034e-11, 4.148866e-11, 4.138473e-11, 4.209266e-11, 
    4.183543e-11, 4.253012e-11, 4.234178e-11, 4.265058e-11, 4.249698e-11, 
    4.24744e-11, 4.22776e-11, 4.215531e-11, 4.184718e-11, 4.159732e-11, 
    4.139974e-11, 4.144563e-11, 4.166282e-11, 4.205765e-11, 4.243294e-11, 
    4.235058e-11, 4.262701e-11, 4.189732e-11, 4.22025e-11, 4.208441e-11, 
    4.239267e-11, 4.171881e-11, 4.22924e-11, 4.157285e-11, 4.163567e-11, 
    4.183032e-11, 4.222332e-11, 4.231049e-11, 4.240371e-11, 4.234616e-11, 
    4.206773e-11, 4.202219e-11, 4.182556e-11, 4.177135e-11, 4.162195e-11, 
    4.149846e-11, 4.161127e-11, 4.172991e-11, 4.206781e-11, 4.237352e-11, 
    4.270813e-11, 4.279021e-11, 4.318331e-11, 4.286318e-11, 4.339213e-11, 
    4.294223e-11, 4.372255e-11, 4.232573e-11, 4.29291e-11, 4.183919e-11, 
    4.19559e-11, 4.216745e-11, 4.26547e-11, 4.239127e-11, 4.269943e-11, 
    4.20204e-11, 4.167034e-11, 4.157999e-11, 4.141174e-11, 4.158383e-11, 
    4.156982e-11, 4.173482e-11, 4.168175e-11, 4.207904e-11, 4.186539e-11, 
    4.247378e-11, 4.269694e-11, 4.333038e-11, 4.372109e-11, 4.412066e-11, 
    4.429766e-11, 4.435161e-11, 4.437416e-11 ;

 F_NIT_vr =
  2.347564e-10, 2.357934e-10, 2.355912e-10, 2.364283e-10, 2.359636e-10, 
    2.365114e-10, 2.349654e-10, 2.35833e-10, 2.352787e-10, 2.348477e-10, 
    2.380524e-10, 2.364637e-10, 2.397047e-10, 2.386894e-10, 2.412401e-10, 
    2.39546e-10, 2.415818e-10, 2.411906e-10, 2.423672e-10, 2.420296e-10, 
    2.435355e-10, 2.425222e-10, 2.443165e-10, 2.43293e-10, 2.434528e-10, 
    2.424876e-10, 2.367849e-10, 2.378563e-10, 2.36721e-10, 2.368738e-10, 
    2.368049e-10, 2.359722e-10, 2.355528e-10, 2.34675e-10, 2.348339e-10, 
    2.354785e-10, 2.369407e-10, 2.364436e-10, 2.376955e-10, 2.376673e-10, 
    2.390624e-10, 2.38433e-10, 2.407807e-10, 2.401126e-10, 2.420434e-10, 
    2.415571e-10, 2.420201e-10, 2.418793e-10, 2.420212e-10, 2.413087e-10, 
    2.416134e-10, 2.409866e-10, 2.385537e-10, 2.392694e-10, 2.371349e-10, 
    2.35853e-10, 2.350024e-10, 2.343994e-10, 2.344842e-10, 2.346467e-10, 
    2.354818e-10, 2.362674e-10, 2.368667e-10, 2.372675e-10, 2.376625e-10, 
    2.388602e-10, 2.394942e-10, 2.409153e-10, 2.406585e-10, 2.41093e-10, 
    2.415085e-10, 2.422062e-10, 2.420912e-10, 2.423984e-10, 2.410802e-10, 
    2.41956e-10, 2.405103e-10, 2.409054e-10, 2.377725e-10, 2.365787e-10, 
    2.360718e-10, 2.356279e-10, 2.345495e-10, 2.35294e-10, 2.350002e-10, 
    2.356982e-10, 2.361421e-10, 2.359221e-10, 2.372782e-10, 2.367503e-10, 
    2.395314e-10, 2.383326e-10, 2.414603e-10, 2.407106e-10, 2.416393e-10, 
    2.411652e-10, 2.419772e-10, 2.41246e-10, 2.425124e-10, 2.427885e-10, 
    2.425994e-10, 2.433242e-10, 2.41204e-10, 2.420177e-10, 2.359173e-10, 
    2.359532e-10, 2.361198e-10, 2.353861e-10, 2.353411e-10, 2.346691e-10, 
    2.352664e-10, 2.35521e-10, 2.361672e-10, 2.365494e-10, 2.369129e-10, 
    2.377133e-10, 2.386074e-10, 2.398589e-10, 2.407589e-10, 2.413624e-10, 
    2.40992e-10, 2.413185e-10, 2.40953e-10, 2.407813e-10, 2.426844e-10, 
    2.416153e-10, 2.432193e-10, 2.431305e-10, 2.424038e-10, 2.431398e-10, 
    2.359779e-10, 2.357714e-10, 2.350561e-10, 2.356154e-10, 2.345956e-10, 
    2.351662e-10, 2.354941e-10, 2.367611e-10, 2.370394e-10, 2.372978e-10, 
    2.378081e-10, 2.384633e-10, 2.396142e-10, 2.40616e-10, 2.415317e-10, 
    2.414642e-10, 2.414877e-10, 2.41692e-10, 2.41185e-10, 2.417748e-10, 
    2.418735e-10, 2.416145e-10, 2.431179e-10, 2.426881e-10, 2.431276e-10, 
    2.428474e-10, 2.358382e-10, 2.361846e-10, 2.359969e-10, 2.363494e-10, 
    2.361005e-10, 2.372052e-10, 2.375363e-10, 2.390879e-10, 2.384504e-10, 
    2.394647e-10, 2.385529e-10, 2.387144e-10, 2.39497e-10, 2.386015e-10, 
    2.4056e-10, 2.392314e-10, 2.416997e-10, 2.403717e-10, 2.417825e-10, 
    2.415257e-10, 2.419498e-10, 2.423302e-10, 2.428082e-10, 2.436917e-10, 
    2.434865e-10, 2.442258e-10, 2.367016e-10, 2.371514e-10, 2.371117e-10, 
    2.375827e-10, 2.379311e-10, 2.386873e-10, 2.399007e-10, 2.394438e-10, 
    2.402818e-10, 2.404503e-10, 2.391761e-10, 2.39958e-10, 2.374504e-10, 
    2.378547e-10, 2.376137e-10, 2.367334e-10, 2.39547e-10, 2.381018e-10, 
    2.407709e-10, 2.399869e-10, 2.422753e-10, 2.411365e-10, 2.433737e-10, 
    2.443316e-10, 2.452334e-10, 2.46288e-10, 2.37397e-10, 2.370906e-10, 
    2.376382e-10, 2.383969e-10, 2.391006e-10, 2.400376e-10, 2.401332e-10, 
    2.403085e-10, 2.40763e-10, 2.411459e-10, 2.403634e-10, 2.412411e-10, 
    2.379484e-10, 2.396724e-10, 2.369717e-10, 2.377843e-10, 2.383488e-10, 
    2.381009e-10, 2.393885e-10, 2.396918e-10, 2.409265e-10, 2.402881e-10, 
    2.440944e-10, 2.424087e-10, 2.470914e-10, 2.45781e-10, 2.369834e-10, 
    2.373949e-10, 2.388291e-10, 2.381464e-10, 2.400995e-10, 2.405808e-10, 
    2.409717e-10, 2.414724e-10, 2.415259e-10, 2.418227e-10, 2.41336e-10, 
    2.41803e-10, 2.40037e-10, 2.408256e-10, 2.386624e-10, 2.391881e-10, 
    2.389459e-10, 2.386801e-10, 2.394993e-10, 2.40373e-10, 2.403914e-10, 
    2.406711e-10, 2.414612e-10, 2.401029e-10, 2.443113e-10, 2.417101e-10, 
    2.378439e-10, 2.386375e-10, 2.387507e-10, 2.38443e-10, 2.40532e-10, 
    2.397745e-10, 2.418155e-10, 2.41263e-10, 2.421674e-10, 2.417178e-10, 
    2.416511e-10, 2.41074e-10, 2.407142e-10, 2.398073e-10, 2.390693e-10, 
    2.384848e-10, 2.386202e-10, 2.392624e-10, 2.404258e-10, 2.415279e-10, 
    2.41286e-10, 2.420956e-10, 2.399528e-10, 2.408507e-10, 2.405031e-10, 
    2.414084e-10, 2.394306e-10, 2.41119e-10, 2.389992e-10, 2.391845e-10, 
    2.397588e-10, 2.409153e-10, 2.411708e-10, 2.414443e-10, 2.41275e-10, 
    2.404571e-10, 2.403228e-10, 2.397432e-10, 2.39583e-10, 2.391419e-10, 
    2.387763e-10, 2.391099e-10, 2.394598e-10, 2.404556e-10, 2.413531e-10, 
    2.423326e-10, 2.425724e-10, 2.43718e-10, 2.42785e-10, 2.443246e-10, 
    2.430151e-10, 2.452822e-10, 2.412162e-10, 2.429815e-10, 2.39785e-10, 
    2.401285e-10, 2.407507e-10, 2.421789e-10, 2.414071e-10, 2.423095e-10, 
    2.403174e-10, 2.392849e-10, 2.390177e-10, 2.3852e-10, 2.390286e-10, 
    2.389873e-10, 2.394744e-10, 2.393173e-10, 2.404879e-10, 2.398589e-10, 
    2.416463e-10, 2.422995e-10, 2.441455e-10, 2.452783e-10, 2.464327e-10, 
    2.469423e-10, 2.470975e-10, 2.471621e-10,
  1.335097e-10, 1.345181e-10, 1.343218e-10, 1.351368e-10, 1.346845e-10, 
    1.352185e-10, 1.337139e-10, 1.345582e-10, 1.34019e-10, 1.336004e-10, 
    1.367235e-10, 1.351732e-10, 1.383408e-10, 1.37347e-10, 1.398483e-10, 
    1.381859e-10, 1.401844e-10, 1.398003e-10, 1.409575e-10, 1.406256e-10, 
    1.421095e-10, 1.411108e-10, 1.428809e-10, 1.418708e-10, 1.420286e-10, 
    1.410779e-10, 1.354847e-10, 1.365301e-10, 1.354229e-10, 1.355717e-10, 
    1.355049e-10, 1.346939e-10, 1.342858e-10, 1.334327e-10, 1.335875e-10, 
    1.342141e-10, 1.356387e-10, 1.351545e-10, 1.363761e-10, 1.363484e-10, 
    1.37713e-10, 1.370971e-10, 1.39398e-10, 1.387427e-10, 1.406395e-10, 
    1.401616e-10, 1.40617e-10, 1.404789e-10, 1.406188e-10, 1.399181e-10, 
    1.402182e-10, 1.396022e-10, 1.372124e-10, 1.379132e-10, 1.358269e-10, 
    1.34578e-10, 1.337509e-10, 1.331651e-10, 1.332479e-10, 1.334057e-10, 
    1.342177e-10, 1.34983e-10, 1.355672e-10, 1.359585e-10, 1.363445e-10, 
    1.375151e-10, 1.381362e-10, 1.395306e-10, 1.392786e-10, 1.397056e-10, 
    1.40114e-10, 1.408007e-10, 1.406876e-10, 1.409904e-10, 1.396944e-10, 
    1.405552e-10, 1.391352e-10, 1.39523e-10, 1.364493e-10, 1.352851e-10, 
    1.347912e-10, 1.343596e-10, 1.333115e-10, 1.340349e-10, 1.337496e-10, 
    1.344289e-10, 1.348612e-10, 1.346473e-10, 1.359692e-10, 1.354547e-10, 
    1.381731e-10, 1.369998e-10, 1.400664e-10, 1.393303e-10, 1.40243e-10, 
    1.39777e-10, 1.405758e-10, 1.398568e-10, 1.411031e-10, 1.41375e-10, 
    1.411892e-10, 1.419035e-10, 1.39817e-10, 1.40617e-10, 1.346413e-10, 
    1.346762e-10, 1.348387e-10, 1.341249e-10, 1.340813e-10, 1.334285e-10, 
    1.340093e-10, 1.342569e-10, 1.348862e-10, 1.35259e-10, 1.356137e-10, 
    1.363947e-10, 1.37269e-10, 1.384949e-10, 1.39378e-10, 1.399711e-10, 
    1.396073e-10, 1.399285e-10, 1.395695e-10, 1.394013e-10, 1.412731e-10, 
    1.40221e-10, 1.418007e-10, 1.417131e-10, 1.409976e-10, 1.41723e-10, 
    1.347007e-10, 1.345e-10, 1.338043e-10, 1.343486e-10, 1.333575e-10, 
    1.339119e-10, 1.342311e-10, 1.354654e-10, 1.357372e-10, 1.359893e-10, 
    1.364879e-10, 1.371286e-10, 1.382553e-10, 1.392382e-10, 1.401378e-10, 
    1.400719e-10, 1.400951e-10, 1.402963e-10, 1.39798e-10, 1.403782e-10, 
    1.404756e-10, 1.402209e-10, 1.417014e-10, 1.412779e-10, 1.417113e-10, 
    1.414354e-10, 1.345652e-10, 1.349029e-10, 1.347204e-10, 1.350637e-10, 
    1.348218e-10, 1.358986e-10, 1.362221e-10, 1.377394e-10, 1.37116e-10, 
    1.381087e-10, 1.372167e-10, 1.373746e-10, 1.381411e-10, 1.372649e-10, 
    1.39184e-10, 1.378818e-10, 1.403041e-10, 1.389999e-10, 1.40386e-10, 
    1.401339e-10, 1.405513e-10, 1.409255e-10, 1.413968e-10, 1.422679e-10, 
    1.42066e-10, 1.427956e-10, 1.35407e-10, 1.358461e-10, 1.358074e-10, 
    1.362675e-10, 1.36608e-10, 1.373473e-10, 1.38536e-10, 1.380886e-10, 
    1.389104e-10, 1.390756e-10, 1.378272e-10, 1.385932e-10, 1.361402e-10, 
    1.365354e-10, 1.363001e-10, 1.354416e-10, 1.381916e-10, 1.367778e-10, 
    1.393926e-10, 1.386237e-10, 1.408722e-10, 1.397523e-10, 1.419549e-10, 
    1.429002e-10, 1.43792e-10, 1.448365e-10, 1.36086e-10, 1.357874e-10, 
    1.363222e-10, 1.370634e-10, 1.377525e-10, 1.386705e-10, 1.387646e-10, 
    1.389368e-10, 1.393834e-10, 1.397593e-10, 1.389913e-10, 1.398536e-10, 
    1.366271e-10, 1.383146e-10, 1.356745e-10, 1.364675e-10, 1.370197e-10, 
    1.367774e-10, 1.380375e-10, 1.383351e-10, 1.395467e-10, 1.389199e-10, 
    1.426667e-10, 1.410046e-10, 1.456336e-10, 1.443347e-10, 1.356831e-10, 
    1.360849e-10, 1.374869e-10, 1.368192e-10, 1.387319e-10, 1.392041e-10, 
    1.395885e-10, 1.400804e-10, 1.401335e-10, 1.404253e-10, 1.399473e-10, 
    1.404064e-10, 1.386725e-10, 1.394464e-10, 1.373264e-10, 1.378413e-10, 
    1.376043e-10, 1.373446e-10, 1.381469e-10, 1.390034e-10, 1.390217e-10, 
    1.392968e-10, 1.400729e-10, 1.387397e-10, 1.428816e-10, 1.403184e-10, 
    1.365236e-10, 1.372998e-10, 1.374108e-10, 1.371099e-10, 1.391568e-10, 
    1.384138e-10, 1.404182e-10, 1.398754e-10, 1.407651e-10, 1.403228e-10, 
    1.402577e-10, 1.396904e-10, 1.393377e-10, 1.384479e-10, 1.377254e-10, 
    1.371535e-10, 1.372864e-10, 1.379149e-10, 1.390559e-10, 1.401383e-10, 
    1.399009e-10, 1.406974e-10, 1.385929e-10, 1.394739e-10, 1.391332e-10, 
    1.400224e-10, 1.380767e-10, 1.397328e-10, 1.376545e-10, 1.378363e-10, 
    1.383991e-10, 1.395337e-10, 1.397853e-10, 1.40054e-10, 1.398882e-10, 
    1.390849e-10, 1.389534e-10, 1.383854e-10, 1.382287e-10, 1.377967e-10, 
    1.374394e-10, 1.377658e-10, 1.38109e-10, 1.390852e-10, 1.399671e-10, 
    1.409309e-10, 1.411671e-10, 1.422968e-10, 1.413769e-10, 1.428959e-10, 
    1.41604e-10, 1.438431e-10, 1.39829e-10, 1.415662e-10, 1.384247e-10, 
    1.38762e-10, 1.393726e-10, 1.407769e-10, 1.400182e-10, 1.409057e-10, 
    1.389483e-10, 1.379366e-10, 1.376753e-10, 1.371882e-10, 1.376864e-10, 
    1.376459e-10, 1.381232e-10, 1.379698e-10, 1.391177e-10, 1.385006e-10, 
    1.402561e-10, 1.408987e-10, 1.42719e-10, 1.43839e-10, 1.449823e-10, 
    1.45488e-10, 1.456421e-10, 1.457065e-10,
  1.248478e-10, 1.259514e-10, 1.257365e-10, 1.26629e-10, 1.261336e-10, 
    1.267185e-10, 1.250712e-10, 1.259953e-10, 1.25405e-10, 1.24947e-10, 
    1.283686e-10, 1.266689e-10, 1.301443e-10, 1.290529e-10, 1.31802e-10, 
    1.299742e-10, 1.321718e-10, 1.317491e-10, 1.330231e-10, 1.326576e-10, 
    1.342925e-10, 1.331919e-10, 1.351434e-10, 1.340294e-10, 1.342034e-10, 
    1.331557e-10, 1.270102e-10, 1.281564e-10, 1.269424e-10, 1.271056e-10, 
    1.270324e-10, 1.261438e-10, 1.25697e-10, 1.247636e-10, 1.249329e-10, 
    1.256186e-10, 1.27179e-10, 1.266484e-10, 1.279875e-10, 1.279572e-10, 
    1.294547e-10, 1.287786e-10, 1.313066e-10, 1.30586e-10, 1.326728e-10, 
    1.321467e-10, 1.326481e-10, 1.32496e-10, 1.326501e-10, 1.318788e-10, 
    1.32209e-10, 1.315312e-10, 1.289051e-10, 1.296746e-10, 1.273853e-10, 
    1.260169e-10, 1.251117e-10, 1.244709e-10, 1.245614e-10, 1.24734e-10, 
    1.256226e-10, 1.264605e-10, 1.271006e-10, 1.275296e-10, 1.279528e-10, 
    1.292374e-10, 1.299196e-10, 1.314525e-10, 1.311753e-10, 1.31645e-10, 
    1.320944e-10, 1.328503e-10, 1.327258e-10, 1.330593e-10, 1.316326e-10, 
    1.325801e-10, 1.310176e-10, 1.314441e-10, 1.280678e-10, 1.267915e-10, 
    1.262505e-10, 1.257778e-10, 1.24631e-10, 1.254225e-10, 1.251102e-10, 
    1.258537e-10, 1.263271e-10, 1.260928e-10, 1.275413e-10, 1.269773e-10, 
    1.299601e-10, 1.286718e-10, 1.32042e-10, 1.312322e-10, 1.322364e-10, 
    1.317236e-10, 1.326027e-10, 1.318114e-10, 1.331835e-10, 1.33483e-10, 
    1.332783e-10, 1.340655e-10, 1.317676e-10, 1.326481e-10, 1.260863e-10, 
    1.261245e-10, 1.263024e-10, 1.255209e-10, 1.254732e-10, 1.24759e-10, 
    1.253944e-10, 1.256654e-10, 1.263545e-10, 1.267629e-10, 1.271516e-10, 
    1.28008e-10, 1.289672e-10, 1.303137e-10, 1.312846e-10, 1.319371e-10, 
    1.315369e-10, 1.318902e-10, 1.314952e-10, 1.313103e-10, 1.333707e-10, 
    1.322121e-10, 1.339521e-10, 1.338556e-10, 1.330672e-10, 1.338665e-10, 
    1.261513e-10, 1.259316e-10, 1.251701e-10, 1.257659e-10, 1.246813e-10, 
    1.252879e-10, 1.256372e-10, 1.269891e-10, 1.27287e-10, 1.275634e-10, 
    1.281101e-10, 1.288132e-10, 1.300504e-10, 1.311309e-10, 1.321206e-10, 
    1.32048e-10, 1.320735e-10, 1.32295e-10, 1.317467e-10, 1.323851e-10, 
    1.324924e-10, 1.32212e-10, 1.338427e-10, 1.33376e-10, 1.338536e-10, 
    1.335496e-10, 1.26003e-10, 1.263728e-10, 1.261729e-10, 1.265489e-10, 
    1.26284e-10, 1.274639e-10, 1.278186e-10, 1.294837e-10, 1.287993e-10, 
    1.298893e-10, 1.289099e-10, 1.290832e-10, 1.299249e-10, 1.289627e-10, 
    1.310712e-10, 1.296401e-10, 1.323036e-10, 1.308688e-10, 1.323937e-10, 
    1.321163e-10, 1.325758e-10, 1.329879e-10, 1.335071e-10, 1.344672e-10, 
    1.342446e-10, 1.350492e-10, 1.26925e-10, 1.274063e-10, 1.273639e-10, 
    1.278683e-10, 1.282419e-10, 1.290532e-10, 1.303589e-10, 1.298672e-10, 
    1.307704e-10, 1.30952e-10, 1.295802e-10, 1.304217e-10, 1.277288e-10, 
    1.281623e-10, 1.279042e-10, 1.26963e-10, 1.299804e-10, 1.284281e-10, 
    1.313007e-10, 1.304552e-10, 1.329291e-10, 1.316963e-10, 1.341222e-10, 
    1.351647e-10, 1.361491e-10, 1.37303e-10, 1.276693e-10, 1.273419e-10, 
    1.279284e-10, 1.287416e-10, 1.294981e-10, 1.305067e-10, 1.306101e-10, 
    1.307995e-10, 1.312906e-10, 1.317041e-10, 1.308594e-10, 1.318078e-10, 
    1.282629e-10, 1.301156e-10, 1.272182e-10, 1.280878e-10, 1.286936e-10, 
    1.284277e-10, 1.298111e-10, 1.301381e-10, 1.314702e-10, 1.307809e-10, 
    1.349071e-10, 1.33075e-10, 1.381844e-10, 1.367485e-10, 1.272276e-10, 
    1.276682e-10, 1.292065e-10, 1.284736e-10, 1.305742e-10, 1.310934e-10, 
    1.315161e-10, 1.320574e-10, 1.321158e-10, 1.32437e-10, 1.319109e-10, 
    1.324162e-10, 1.305089e-10, 1.313598e-10, 1.290303e-10, 1.295956e-10, 
    1.293354e-10, 1.290502e-10, 1.299313e-10, 1.308726e-10, 1.308928e-10, 
    1.311953e-10, 1.320491e-10, 1.305827e-10, 1.351442e-10, 1.323194e-10, 
    1.281493e-10, 1.29001e-10, 1.291229e-10, 1.287926e-10, 1.310413e-10, 
    1.302246e-10, 1.324292e-10, 1.318319e-10, 1.328112e-10, 1.323241e-10, 
    1.322526e-10, 1.316283e-10, 1.312402e-10, 1.30262e-10, 1.294684e-10, 
    1.288405e-10, 1.289863e-10, 1.296765e-10, 1.309303e-10, 1.321211e-10, 
    1.318599e-10, 1.327366e-10, 1.304214e-10, 1.313901e-10, 1.310153e-10, 
    1.319935e-10, 1.298542e-10, 1.316749e-10, 1.293905e-10, 1.295901e-10, 
    1.302084e-10, 1.314559e-10, 1.317326e-10, 1.320283e-10, 1.318458e-10, 
    1.309622e-10, 1.308177e-10, 1.301934e-10, 1.300212e-10, 1.295466e-10, 
    1.291543e-10, 1.295127e-10, 1.298896e-10, 1.309626e-10, 1.319327e-10, 
    1.329937e-10, 1.332539e-10, 1.344991e-10, 1.334851e-10, 1.3516e-10, 
    1.337354e-10, 1.362055e-10, 1.317808e-10, 1.336937e-10, 1.302366e-10, 
    1.306072e-10, 1.312787e-10, 1.328242e-10, 1.319889e-10, 1.32966e-10, 
    1.308121e-10, 1.297003e-10, 1.294133e-10, 1.288786e-10, 1.294256e-10, 
    1.29381e-10, 1.299053e-10, 1.297367e-10, 1.309983e-10, 1.3032e-10, 
    1.322507e-10, 1.329583e-10, 1.349648e-10, 1.36201e-10, 1.374642e-10, 
    1.380233e-10, 1.381937e-10, 1.38265e-10,
  1.280645e-10, 1.292799e-10, 1.290432e-10, 1.300266e-10, 1.294806e-10, 
    1.301252e-10, 1.283105e-10, 1.293282e-10, 1.286781e-10, 1.281737e-10, 
    1.319453e-10, 1.300705e-10, 1.339062e-10, 1.327006e-10, 1.35739e-10, 
    1.337183e-10, 1.361483e-10, 1.356805e-10, 1.370906e-10, 1.366859e-10, 
    1.384971e-10, 1.372776e-10, 1.394404e-10, 1.382054e-10, 1.383982e-10, 
    1.372374e-10, 1.304468e-10, 1.317112e-10, 1.30372e-10, 1.305519e-10, 
    1.304712e-10, 1.294919e-10, 1.289997e-10, 1.279718e-10, 1.281581e-10, 
    1.289132e-10, 1.306329e-10, 1.300479e-10, 1.315246e-10, 1.314911e-10, 
    1.331443e-10, 1.323977e-10, 1.35191e-10, 1.343943e-10, 1.367028e-10, 
    1.361205e-10, 1.366754e-10, 1.36507e-10, 1.366776e-10, 1.35824e-10, 
    1.361894e-10, 1.354395e-10, 1.325374e-10, 1.333872e-10, 1.308604e-10, 
    1.293522e-10, 1.28355e-10, 1.276497e-10, 1.277493e-10, 1.279393e-10, 
    1.289177e-10, 1.298408e-10, 1.305464e-10, 1.310194e-10, 1.314863e-10, 
    1.329044e-10, 1.336579e-10, 1.353524e-10, 1.350458e-10, 1.355654e-10, 
    1.360626e-10, 1.368993e-10, 1.367614e-10, 1.371307e-10, 1.355517e-10, 
    1.366001e-10, 1.348714e-10, 1.353432e-10, 1.316134e-10, 1.302056e-10, 
    1.296094e-10, 1.290886e-10, 1.278259e-10, 1.286973e-10, 1.283534e-10, 
    1.291722e-10, 1.296937e-10, 1.294357e-10, 1.310324e-10, 1.304105e-10, 
    1.337026e-10, 1.322798e-10, 1.360046e-10, 1.351087e-10, 1.362197e-10, 
    1.356523e-10, 1.366252e-10, 1.357494e-10, 1.372682e-10, 1.376e-10, 
    1.373733e-10, 1.382454e-10, 1.357009e-10, 1.366754e-10, 1.294284e-10, 
    1.294705e-10, 1.296666e-10, 1.288057e-10, 1.287531e-10, 1.279667e-10, 
    1.286663e-10, 1.289648e-10, 1.29724e-10, 1.301741e-10, 1.306026e-10, 
    1.315472e-10, 1.32606e-10, 1.340933e-10, 1.351667e-10, 1.358886e-10, 
    1.354457e-10, 1.358366e-10, 1.353997e-10, 1.351951e-10, 1.374757e-10, 
    1.361928e-10, 1.381198e-10, 1.380128e-10, 1.371395e-10, 1.380248e-10, 
    1.295001e-10, 1.29258e-10, 1.284193e-10, 1.290754e-10, 1.278812e-10, 
    1.28549e-10, 1.289338e-10, 1.304235e-10, 1.307519e-10, 1.310568e-10, 
    1.316599e-10, 1.324359e-10, 1.338023e-10, 1.349968e-10, 1.360915e-10, 
    1.360112e-10, 1.360395e-10, 1.362846e-10, 1.356778e-10, 1.363843e-10, 
    1.365031e-10, 1.361927e-10, 1.379985e-10, 1.374814e-10, 1.380105e-10, 
    1.376737e-10, 1.293367e-10, 1.297442e-10, 1.295239e-10, 1.299383e-10, 
    1.296463e-10, 1.309471e-10, 1.313384e-10, 1.331764e-10, 1.324206e-10, 
    1.336244e-10, 1.325426e-10, 1.32734e-10, 1.336638e-10, 1.32601e-10, 
    1.349308e-10, 1.333491e-10, 1.362941e-10, 1.347071e-10, 1.363939e-10, 
    1.360868e-10, 1.365954e-10, 1.370516e-10, 1.376266e-10, 1.386907e-10, 
    1.384439e-10, 1.39336e-10, 1.303529e-10, 1.308836e-10, 1.308368e-10, 
    1.313931e-10, 1.318053e-10, 1.327009e-10, 1.341432e-10, 1.336e-10, 
    1.345981e-10, 1.347989e-10, 1.332828e-10, 1.342127e-10, 1.312393e-10, 
    1.317175e-10, 1.314327e-10, 1.303947e-10, 1.337251e-10, 1.320109e-10, 
    1.351845e-10, 1.342497e-10, 1.369865e-10, 1.356222e-10, 1.383082e-10, 
    1.394641e-10, 1.405562e-10, 1.418376e-10, 1.311736e-10, 1.308125e-10, 
    1.314594e-10, 1.323569e-10, 1.331922e-10, 1.343066e-10, 1.344209e-10, 
    1.346303e-10, 1.351733e-10, 1.356307e-10, 1.346965e-10, 1.357454e-10, 
    1.318286e-10, 1.338744e-10, 1.306761e-10, 1.316353e-10, 1.323039e-10, 
    1.320104e-10, 1.335379e-10, 1.338992e-10, 1.35372e-10, 1.346097e-10, 
    1.391784e-10, 1.371481e-10, 1.428169e-10, 1.412217e-10, 1.306865e-10, 
    1.311724e-10, 1.328701e-10, 1.32061e-10, 1.343812e-10, 1.349553e-10, 
    1.354228e-10, 1.360216e-10, 1.360863e-10, 1.364418e-10, 1.358595e-10, 
    1.364187e-10, 1.34309e-10, 1.352499e-10, 1.326755e-10, 1.332999e-10, 
    1.330125e-10, 1.326976e-10, 1.336707e-10, 1.347112e-10, 1.347334e-10, 
    1.350679e-10, 1.360127e-10, 1.343906e-10, 1.394415e-10, 1.363118e-10, 
    1.317032e-10, 1.326433e-10, 1.327778e-10, 1.324131e-10, 1.348977e-10, 
    1.339949e-10, 1.364331e-10, 1.35772e-10, 1.368559e-10, 1.363168e-10, 
    1.362376e-10, 1.355469e-10, 1.351177e-10, 1.340362e-10, 1.331593e-10, 
    1.32466e-10, 1.32627e-10, 1.333892e-10, 1.34775e-10, 1.360922e-10, 
    1.358031e-10, 1.367734e-10, 1.342123e-10, 1.352834e-10, 1.34869e-10, 
    1.359509e-10, 1.335855e-10, 1.355986e-10, 1.330733e-10, 1.332938e-10, 
    1.33977e-10, 1.353562e-10, 1.356623e-10, 1.359894e-10, 1.357875e-10, 
    1.348102e-10, 1.346504e-10, 1.339603e-10, 1.337701e-10, 1.332458e-10, 
    1.328124e-10, 1.332083e-10, 1.336247e-10, 1.348106e-10, 1.358836e-10, 
    1.370581e-10, 1.373463e-10, 1.387261e-10, 1.376024e-10, 1.394591e-10, 
    1.378798e-10, 1.40619e-10, 1.357157e-10, 1.378335e-10, 1.340081e-10, 
    1.344177e-10, 1.351602e-10, 1.368704e-10, 1.359458e-10, 1.370274e-10, 
    1.346442e-10, 1.334156e-10, 1.330986e-10, 1.325081e-10, 1.331121e-10, 
    1.330629e-10, 1.33642e-10, 1.334558e-10, 1.348501e-10, 1.341003e-10, 
    1.362356e-10, 1.370189e-10, 1.392424e-10, 1.406139e-10, 1.420165e-10, 
    1.426379e-10, 1.428273e-10, 1.429065e-10,
  1.381445e-10, 1.394321e-10, 1.391812e-10, 1.402237e-10, 1.396448e-10, 
    1.403282e-10, 1.38405e-10, 1.394834e-10, 1.387944e-10, 1.382601e-10, 
    1.422596e-10, 1.402703e-10, 1.443425e-10, 1.430614e-10, 1.462921e-10, 
    1.441428e-10, 1.467276e-10, 1.462297e-10, 1.477311e-10, 1.473001e-10, 
    1.492303e-10, 1.479303e-10, 1.502365e-10, 1.489192e-10, 1.491249e-10, 
    1.478875e-10, 1.406692e-10, 1.420111e-10, 1.4059e-10, 1.407808e-10, 
    1.406951e-10, 1.396568e-10, 1.391352e-10, 1.380463e-10, 1.382436e-10, 
    1.390436e-10, 1.408667e-10, 1.402462e-10, 1.418127e-10, 1.417772e-10, 
    1.435327e-10, 1.427397e-10, 1.457088e-10, 1.448613e-10, 1.47318e-10, 
    1.46698e-10, 1.472889e-10, 1.471096e-10, 1.472912e-10, 1.463824e-10, 
    1.467714e-10, 1.459732e-10, 1.42888e-10, 1.437908e-10, 1.411079e-10, 
    1.395088e-10, 1.384522e-10, 1.377052e-10, 1.378107e-10, 1.380119e-10, 
    1.390482e-10, 1.400266e-10, 1.407749e-10, 1.412767e-10, 1.417721e-10, 
    1.432781e-10, 1.440786e-10, 1.458806e-10, 1.455543e-10, 1.461072e-10, 
    1.466364e-10, 1.475274e-10, 1.473805e-10, 1.477739e-10, 1.460925e-10, 
    1.472087e-10, 1.453687e-10, 1.458707e-10, 1.419073e-10, 1.404134e-10, 
    1.397815e-10, 1.392294e-10, 1.378918e-10, 1.388148e-10, 1.384505e-10, 
    1.393179e-10, 1.398708e-10, 1.395972e-10, 1.412904e-10, 1.406308e-10, 
    1.441261e-10, 1.426145e-10, 1.465746e-10, 1.456213e-10, 1.468036e-10, 
    1.461996e-10, 1.472355e-10, 1.46303e-10, 1.479204e-10, 1.48274e-10, 
    1.480323e-10, 1.489618e-10, 1.462514e-10, 1.472889e-10, 1.395895e-10, 
    1.396341e-10, 1.39842e-10, 1.389296e-10, 1.388739e-10, 1.380409e-10, 
    1.387819e-10, 1.390982e-10, 1.399028e-10, 1.4038e-10, 1.408345e-10, 
    1.418368e-10, 1.429609e-10, 1.445414e-10, 1.45683e-10, 1.464511e-10, 
    1.459798e-10, 1.463958e-10, 1.459308e-10, 1.457131e-10, 1.481414e-10, 
    1.467751e-10, 1.488279e-10, 1.487138e-10, 1.477832e-10, 1.487267e-10, 
    1.396654e-10, 1.394089e-10, 1.385203e-10, 1.392154e-10, 1.379504e-10, 
    1.386577e-10, 1.390654e-10, 1.406446e-10, 1.409929e-10, 1.413163e-10, 
    1.419564e-10, 1.427802e-10, 1.442321e-10, 1.455022e-10, 1.466672e-10, 
    1.465816e-10, 1.466118e-10, 1.468727e-10, 1.462268e-10, 1.469789e-10, 
    1.471054e-10, 1.467749e-10, 1.486986e-10, 1.481475e-10, 1.487114e-10, 
    1.483525e-10, 1.394922e-10, 1.399242e-10, 1.396907e-10, 1.4013e-10, 
    1.398205e-10, 1.412001e-10, 1.416152e-10, 1.435669e-10, 1.42764e-10, 
    1.44043e-10, 1.428936e-10, 1.430969e-10, 1.44085e-10, 1.429556e-10, 
    1.454321e-10, 1.437505e-10, 1.468829e-10, 1.451941e-10, 1.469891e-10, 
    1.466621e-10, 1.472036e-10, 1.476896e-10, 1.483023e-10, 1.494367e-10, 
    1.491735e-10, 1.50125e-10, 1.405696e-10, 1.411326e-10, 1.410829e-10, 
    1.416733e-10, 1.421108e-10, 1.430617e-10, 1.445945e-10, 1.44017e-10, 
    1.450781e-10, 1.452917e-10, 1.436799e-10, 1.446684e-10, 1.4151e-10, 
    1.420176e-10, 1.417152e-10, 1.40614e-10, 1.4415e-10, 1.423291e-10, 
    1.457019e-10, 1.447076e-10, 1.476203e-10, 1.461676e-10, 1.490288e-10, 
    1.502619e-10, 1.514275e-10, 1.527967e-10, 1.414403e-10, 1.410572e-10, 
    1.417435e-10, 1.426964e-10, 1.435837e-10, 1.447682e-10, 1.448897e-10, 
    1.451123e-10, 1.456899e-10, 1.461766e-10, 1.451828e-10, 1.462988e-10, 
    1.421357e-10, 1.443086e-10, 1.409125e-10, 1.419304e-10, 1.426401e-10, 
    1.423285e-10, 1.43951e-10, 1.44335e-10, 1.459014e-10, 1.450904e-10, 
    1.499571e-10, 1.477925e-10, 1.538438e-10, 1.521385e-10, 1.409235e-10, 
    1.414389e-10, 1.432415e-10, 1.423822e-10, 1.448474e-10, 1.45458e-10, 
    1.459554e-10, 1.465927e-10, 1.466616e-10, 1.470401e-10, 1.464202e-10, 
    1.470155e-10, 1.447707e-10, 1.457714e-10, 1.430348e-10, 1.436981e-10, 
    1.433927e-10, 1.430582e-10, 1.440921e-10, 1.451985e-10, 1.452221e-10, 
    1.455779e-10, 1.465835e-10, 1.448575e-10, 1.50238e-10, 1.469019e-10, 
    1.420023e-10, 1.430007e-10, 1.431435e-10, 1.42756e-10, 1.453967e-10, 
    1.444367e-10, 1.470308e-10, 1.463271e-10, 1.474812e-10, 1.46907e-10, 
    1.468227e-10, 1.460874e-10, 1.456308e-10, 1.444807e-10, 1.435488e-10, 
    1.428122e-10, 1.429833e-10, 1.43793e-10, 1.452663e-10, 1.466679e-10, 
    1.463602e-10, 1.473933e-10, 1.446679e-10, 1.458072e-10, 1.453662e-10, 
    1.465175e-10, 1.440016e-10, 1.461428e-10, 1.434573e-10, 1.436916e-10, 
    1.444177e-10, 1.458847e-10, 1.462103e-10, 1.465585e-10, 1.463435e-10, 
    1.453038e-10, 1.451338e-10, 1.444e-10, 1.441978e-10, 1.436406e-10, 
    1.431802e-10, 1.436008e-10, 1.440433e-10, 1.453042e-10, 1.464459e-10, 
    1.476965e-10, 1.480035e-10, 1.494746e-10, 1.482766e-10, 1.502567e-10, 
    1.485725e-10, 1.514948e-10, 1.462672e-10, 1.485229e-10, 1.444507e-10, 
    1.448863e-10, 1.456761e-10, 1.474967e-10, 1.465121e-10, 1.476639e-10, 
    1.451271e-10, 1.438211e-10, 1.434841e-10, 1.428569e-10, 1.434985e-10, 
    1.434462e-10, 1.440616e-10, 1.438637e-10, 1.453461e-10, 1.445487e-10, 
    1.468206e-10, 1.476548e-10, 1.500252e-10, 1.514892e-10, 1.529879e-10, 
    1.536523e-10, 1.538548e-10, 1.539396e-10,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GC_HEAT1 =
  24532.13, 24552.02, 24548.12, 24564.4, 24555.33, 24566.04, 24536.13, 
    24552.81, 24542.13, 24533.9, 24596.72, 24565.13, 24630.54, 24609.63, 
    24662.6, 24627.26, 24669.87, 24661.57, 24686.78, 24679.49, 24712.5, 
    24690.16, 24730.1, 24707.11, 24710.67, 24689.44, 24571.42, 24592.75, 
    24570.17, 24573.18, 24571.83, 24555.52, 24547.4, 24530.63, 24533.65, 
    24545.98, 24574.54, 24564.75, 24589.58, 24589.02, 24617.28, 24604.44, 
    24652.95, 24639.05, 24679.79, 24669.37, 24679.3, 24676.28, 24679.34, 
    24664.11, 24670.6, 24657.31, 24606.83, 24621.49, 24578.37, 24553.21, 
    24536.86, 24525.42, 24527.03, 24530.1, 24546.06, 24561.3, 24573.09, 
    24581.05, 24588.94, 24613.14, 24626.2, 24655.78, 24650.4, 24659.53, 
    24668.34, 24683.33, 24680.85, 24687.51, 24659.29, 24677.95, 24647.35, 
    24655.62, 24591.09, 24567.38, 24557.47, 24548.87, 24528.26, 24542.45, 
    24536.83, 24550.24, 24558.86, 24554.59, 24581.27, 24570.81, 24626.98, 
    24602.42, 24667.31, 24651.5, 24671.14, 24661.07, 24678.4, 24662.79, 
    24690, 24696.03, 24691.9, 24707.85, 24661.93, 24679.3, 24554.47, 
    24555.16, 24558.41, 24544.22, 24543.36, 24530.54, 24541.94, 24546.83, 
    24559.36, 24566.86, 24574.03, 24589.96, 24608.01, 24633.82, 24652.52, 
    24665.25, 24657.42, 24664.33, 24656.61, 24653.02, 24693.76, 24670.66, 
    24705.54, 24703.57, 24687.67, 24703.79, 24555.65, 24551.65, 24537.9, 
    24548.65, 24529.16, 24540.02, 24546.32, 24571.03, 24576.54, 24581.69, 
    24591.87, 24605.09, 24628.72, 24649.54, 24668.86, 24667.43, 24667.93, 
    24672.3, 24661.52, 24674.08, 24676.21, 24670.66, 24703.31, 24693.87, 
    24703.53, 24697.37, 24552.95, 24559.7, 24556.05, 24562.93, 24558.07, 
    24579.83, 24586.44, 24617.84, 24604.83, 24625.62, 24606.92, 24610.21, 
    24626.31, 24607.92, 24648.39, 24620.83, 24672.47, 24644.49, 24674.25, 
    24668.77, 24677.86, 24686.08, 24696.51, 24716.09, 24711.51, 24728.13, 
    24569.84, 24578.76, 24577.97, 24587.36, 24594.34, 24609.63, 24634.7, 
    24625.19, 24642.59, 24646.09, 24619.68, 24635.91, 24584.77, 24592.85, 
    24588.03, 24570.54, 24627.38, 24597.83, 24652.83, 24636.55, 24684.9, 
    24660.54, 24709.01, 24730.55, 24751.25, 24775.9, 24583.66, 24577.56, 
    24588.48, 24603.74, 24618.11, 24637.54, 24639.51, 24643.15, 24652.63, 
    24660.69, 24644.3, 24662.71, 24594.74, 24629.98, 24575.27, 24591.46, 
    24602.83, 24597.82, 24624.11, 24630.42, 24656.12, 24642.79, 24725.18, 
    24687.82, 24794.88, 24764.07, 24575.44, 24583.64, 24612.55, 24598.69, 
    24638.83, 24648.82, 24657.02, 24667.62, 24668.77, 24675.11, 24664.74, 
    24674.7, 24637.58, 24653.98, 24609.2, 24619.98, 24615, 24609.58, 
    24626.42, 24644.56, 24644.95, 24650.79, 24667.46, 24638.99, 24730.12, 
    24672.79, 24592.61, 24608.65, 24610.96, 24604.7, 24647.81, 24632.09, 
    24674.96, 24663.19, 24682.55, 24672.88, 24671.46, 24659.21, 24651.66, 
    24632.82, 24617.54, 24605.6, 24608.37, 24621.53, 24645.67, 24668.87, 
    24663.74, 24681.06, 24635.9, 24654.57, 24647.31, 24666.36, 24624.94, 
    24660.12, 24616.05, 24619.87, 24631.78, 24655.85, 24661.24, 24667.04, 
    24663.46, 24646.29, 24643.5, 24631.49, 24628.16, 24619.04, 24611.55, 
    24618.39, 24625.62, 24646.29, 24665.16, 24686.2, 24691.41, 24716.75, 
    24696.07, 24730.46, 24701.14, 24752.45, 24662.19, 24700.29, 24632.32, 
    24639.46, 24652.41, 24682.81, 24666.27, 24685.64, 24643.39, 24621.99, 
    24616.49, 24606.33, 24616.72, 24615.88, 24625.92, 24622.68, 24646.98, 
    24633.94, 24671.43, 24685.49, 24726.38, 24752.35, 24779.35, 24791.39, 
    24795.08, 24796.63 ;

 GC_ICE1 =
  17606.22, 17637.98, 17631.75, 17657.75, 17643.27, 17660.38, 17612.6, 
    17639.26, 17622.19, 17609.05, 17709.36, 17658.92, 17763.31, 17729.95, 
    17814.36, 17758.07, 17825.92, 17812.71, 17852.83, 17841.22, 17893.74, 
    17858.21, 17921.73, 17885.17, 17890.83, 17857.05, 17668.96, 17703.02, 
    17666.97, 17671.78, 17669.62, 17643.57, 17630.62, 17603.81, 17608.65, 
    17628.34, 17673.96, 17658.32, 17697.96, 17697.06, 17742.16, 17721.66, 
    17798.98, 17776.87, 17841.71, 17825.13, 17840.92, 17836.12, 17840.99, 
    17816.75, 17827.08, 17805.94, 17725.48, 17748.88, 17680.07, 17639.89, 
    17613.76, 17595.49, 17598.06, 17602.97, 17628.46, 17652.81, 17671.63, 
    17684.36, 17696.93, 17735.56, 17756.39, 17803.5, 17794.93, 17809.47, 
    17823.49, 17847.34, 17843.39, 17853.98, 17809.08, 17838.77, 17790.08, 
    17803.24, 17700.38, 17662.52, 17646.68, 17632.95, 17600.04, 17622.69, 
    17613.72, 17635.14, 17648.91, 17642.09, 17684.71, 17667.99, 17757.63, 
    17718.45, 17821.85, 17796.69, 17827.94, 17811.91, 17839.49, 17814.64, 
    17857.94, 17867.53, 17860.97, 17886.34, 17813.28, 17840.93, 17641.9, 
    17643.01, 17648.19, 17625.53, 17624.15, 17603.68, 17621.88, 17629.7, 
    17649.71, 17661.68, 17673.14, 17698.58, 17727.36, 17768.54, 17798.3, 
    17818.57, 17806.11, 17817.1, 17804.82, 17799.1, 17863.93, 17827.18, 
    17882.66, 17879.54, 17854.23, 17879.89, 17643.79, 17637.4, 17615.44, 
    17632.6, 17601.47, 17618.82, 17628.88, 17668.34, 17677.15, 17685.36, 
    17701.62, 17722.71, 17760.41, 17793.57, 17824.31, 17822.03, 17822.83, 
    17829.79, 17812.63, 17832.62, 17836, 17827.18, 17879.12, 17864.1, 
    17879.47, 17869.67, 17639.47, 17650.25, 17644.42, 17655.4, 17647.66, 
    17682.41, 17692.95, 17743.05, 17722.29, 17755.46, 17725.62, 17730.87, 
    17756.56, 17727.22, 17791.73, 17747.82, 17830.05, 17785.53, 17832.89, 
    17824.17, 17838.64, 17851.71, 17868.3, 17899.44, 17892.17, 17918.61, 
    17666.45, 17680.69, 17679.43, 17694.42, 17705.56, 17729.96, 17769.94, 
    17754.78, 17782.5, 17788.07, 17745.98, 17771.88, 17690.28, 17703.19, 
    17695.49, 17667.57, 17758.26, 17711.13, 17798.8, 17772.89, 17849.84, 
    17811.07, 17888.18, 17922.44, 17955.35, 17994.51, 17688.52, 17678.78, 
    17696.21, 17720.55, 17743.48, 17774.46, 17777.61, 17783.39, 17798.49, 
    17811.3, 17785.23, 17814.53, 17706.19, 17762.42, 17675.12, 17700.96, 
    17719.11, 17711.12, 17753.05, 17763.11, 17804.04, 17782.82, 17913.91, 
    17854.48, 18024.59, 17975.74, 17675.39, 17688.48, 17734.61, 17712.49, 
    17776.51, 17792.41, 17805.47, 17822.33, 17824.16, 17834.26, 17817.75, 
    17833.6, 17774.53, 17800.63, 17729.27, 17746.46, 17738.53, 17729.87, 
    17756.74, 17785.64, 17786.25, 17795.55, 17822.09, 17776.77, 17921.77, 
    17830.57, 17702.79, 17728.39, 17732.07, 17722.08, 17790.81, 17765.78, 
    17834.01, 17815.28, 17846.09, 17830.7, 17828.45, 17808.95, 17796.94, 
    17766.94, 17742.57, 17723.53, 17727.94, 17748.93, 17787.41, 17824.33, 
    17816.16, 17843.73, 17771.86, 17801.57, 17790.02, 17820.33, 17754.38, 
    17810.41, 17740.2, 17746.29, 17765.28, 17803.61, 17812.19, 17821.42, 
    17815.72, 17788.38, 17783.95, 17764.82, 17759.51, 17744.96, 17733.02, 
    17743.93, 17755.47, 17788.39, 17818.43, 17851.89, 17860.19, 17900.49, 
    17867.61, 17922.3, 17875.67, 17957.27, 17813.7, 17874.32, 17766.15, 
    17777.52, 17798.12, 17846.51, 17820.19, 17851.01, 17783.78, 17749.66, 
    17740.9, 17724.68, 17741.27, 17739.91, 17755.94, 17750.77, 17789.49, 
    17768.73, 17828.39, 17850.77, 17915.81, 17957.11, 17999.98, 18019.06, 
    18024.91, 18027.37 ;

 GC_LIQ1 =
  5232.783, 5234.812, 5234.414, 5236.075, 5235.15, 5236.243, 5233.19, 
    5234.893, 5233.803, 5232.963, 5239.384, 5236.15, 5242.863, 5240.711, 
    5246.213, 5242.525, 5246.975, 5246.105, 5248.749, 5247.983, 5251.45, 
    5249.104, 5253.299, 5250.884, 5251.258, 5249.027, 5236.792, 5238.976, 
    5236.664, 5236.972, 5236.833, 5235.169, 5234.341, 5232.629, 5232.938, 
    5234.196, 5237.111, 5236.111, 5238.65, 5238.592, 5241.499, 5240.177, 
    5245.201, 5243.746, 5248.015, 5246.923, 5247.963, 5247.647, 5247.968, 
    5246.371, 5247.052, 5245.659, 5240.423, 5241.932, 5237.501, 5234.934, 
    5233.265, 5232.098, 5232.262, 5232.576, 5234.204, 5235.759, 5236.962, 
    5237.775, 5238.583, 5241.073, 5242.417, 5245.499, 5244.935, 5245.892, 
    5246.815, 5248.386, 5248.126, 5248.825, 5245.866, 5247.822, 5244.615, 
    5245.481, 5238.805, 5236.38, 5235.368, 5234.49, 5232.388, 5233.835, 
    5233.262, 5234.63, 5235.51, 5235.074, 5237.798, 5236.73, 5242.498, 
    5239.97, 5246.707, 5245.05, 5247.108, 5246.052, 5247.869, 5246.232, 
    5249.086, 5249.719, 5249.286, 5250.961, 5246.143, 5247.964, 5235.062, 
    5235.133, 5235.464, 5234.016, 5233.928, 5232.621, 5233.783, 5234.283, 
    5235.562, 5236.326, 5237.059, 5238.689, 5240.544, 5243.201, 5245.157, 
    5246.491, 5245.67, 5246.395, 5245.585, 5245.208, 5249.481, 5247.058, 
    5250.718, 5250.512, 5248.841, 5250.535, 5235.183, 5234.775, 5233.372, 
    5234.468, 5232.479, 5233.587, 5234.23, 5236.752, 5237.315, 5237.84, 
    5238.886, 5240.245, 5242.676, 5244.845, 5246.869, 5246.719, 5246.772, 
    5247.229, 5246.1, 5247.417, 5247.64, 5247.058, 5250.484, 5249.492, 
    5250.508, 5249.86, 5234.907, 5235.596, 5235.223, 5235.925, 5235.43, 
    5237.651, 5238.327, 5241.556, 5240.217, 5242.357, 5240.433, 5240.771, 
    5242.428, 5240.536, 5244.724, 5241.864, 5247.248, 5244.315, 5247.435, 
    5246.86, 5247.813, 5248.675, 5249.77, 5251.827, 5251.346, 5253.093, 
    5236.631, 5237.542, 5237.461, 5238.422, 5239.139, 5240.712, 5243.291, 
    5242.313, 5244.116, 5244.483, 5241.746, 5243.417, 5238.155, 5238.986, 
    5238.491, 5236.703, 5242.538, 5239.499, 5245.189, 5243.484, 5248.551, 
    5245.997, 5251.083, 5253.346, 5255.528, 5258.146, 5238.042, 5237.419, 
    5238.537, 5240.105, 5241.584, 5243.587, 5243.794, 5244.175, 5245.168, 
    5246.012, 5244.296, 5246.225, 5239.18, 5242.806, 5237.185, 5238.843, 
    5240.012, 5239.498, 5242.202, 5242.851, 5245.535, 5244.137, 5252.783, 
    5248.858, 5260.191, 5256.88, 5237.203, 5238.04, 5241.012, 5239.586, 
    5243.722, 5244.769, 5245.628, 5246.739, 5246.859, 5247.524, 5246.437, 
    5247.481, 5243.591, 5245.31, 5240.667, 5241.776, 5241.265, 5240.706, 
    5242.44, 5244.323, 5244.363, 5244.975, 5246.723, 5243.739, 5253.302, 
    5247.281, 5238.961, 5240.611, 5240.848, 5240.204, 5244.663, 5243.023, 
    5247.508, 5246.274, 5248.304, 5247.29, 5247.142, 5245.857, 5245.066, 
    5243.098, 5241.526, 5240.297, 5240.582, 5241.936, 5244.439, 5246.87, 
    5246.332, 5248.148, 5243.416, 5245.372, 5244.611, 5246.607, 5242.287, 
    5245.954, 5241.373, 5241.765, 5242.991, 5245.506, 5246.071, 5246.679, 
    5246.303, 5244.503, 5244.212, 5242.961, 5242.619, 5241.68, 5240.91, 
    5241.613, 5242.357, 5244.504, 5246.482, 5248.687, 5249.234, 5251.896, 
    5249.724, 5253.337, 5250.257, 5255.655, 5246.17, 5250.167, 5243.047, 
    5243.789, 5245.145, 5248.332, 5246.598, 5248.629, 5244.2, 5241.983, 
    5241.417, 5240.372, 5241.441, 5241.354, 5242.388, 5242.055, 5244.576, 
    5243.213, 5247.138, 5248.613, 5252.908, 5255.645, 5258.517, 5259.814, 
    5260.213, 5260.38 ;

 GPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GROSS_NMIN =
  8.956448e-09, 8.995829e-09, 8.988173e-09, 9.019937e-09, 9.002316e-09, 
    9.023116e-09, 8.964432e-09, 8.997393e-09, 8.976351e-09, 8.959993e-09, 
    9.081578e-09, 9.021353e-09, 9.144131e-09, 9.105723e-09, 9.202203e-09, 
    9.138154e-09, 9.215118e-09, 9.200354e-09, 9.244784e-09, 9.232056e-09, 
    9.288888e-09, 9.250659e-09, 9.318345e-09, 9.279757e-09, 9.285794e-09, 
    9.249399e-09, 9.033473e-09, 9.074081e-09, 9.031067e-09, 9.036857e-09, 
    9.034259e-09, 9.00268e-09, 8.986768e-09, 8.953438e-09, 8.959488e-09, 
    8.983968e-09, 9.039462e-09, 9.020623e-09, 9.068097e-09, 9.067025e-09, 
    9.119877e-09, 9.096047e-09, 9.184878e-09, 9.159631e-09, 9.232587e-09, 
    9.21424e-09, 9.231726e-09, 9.226423e-09, 9.231795e-09, 9.204886e-09, 
    9.216415e-09, 9.192736e-09, 9.100511e-09, 9.127616e-09, 9.046775e-09, 
    8.998167e-09, 8.965878e-09, 8.942965e-09, 8.946205e-09, 8.95238e-09, 
    8.984111e-09, 9.013944e-09, 9.036679e-09, 9.051886e-09, 9.066871e-09, 
    9.112229e-09, 9.136234e-09, 9.189984e-09, 9.180283e-09, 9.196716e-09, 
    9.212415e-09, 9.238772e-09, 9.234433e-09, 9.246046e-09, 9.196282e-09, 
    9.229355e-09, 9.174758e-09, 9.189691e-09, 9.070948e-09, 9.025706e-09, 
    9.006478e-09, 8.989645e-09, 8.948695e-09, 8.976975e-09, 8.965827e-09, 
    8.992347e-09, 9.009199e-09, 9.000864e-09, 9.052303e-09, 9.032305e-09, 
    9.137657e-09, 9.092279e-09, 9.210583e-09, 9.182274e-09, 9.217369e-09, 
    9.199461e-09, 9.230146e-09, 9.202529e-09, 9.250367e-09, 9.260784e-09, 
    9.253665e-09, 9.281009e-09, 9.200998e-09, 9.231726e-09, 9.00063e-09, 
    9.00199e-09, 9.008323e-09, 8.980487e-09, 8.978783e-09, 8.953272e-09, 
    8.975972e-09, 8.985638e-09, 9.010176e-09, 9.02469e-09, 9.038487e-09, 
    9.068823e-09, 9.102703e-09, 9.150076e-09, 9.184109e-09, 9.206922e-09, 
    9.192934e-09, 9.205284e-09, 9.191478e-09, 9.185007e-09, 9.256881e-09, 
    9.216523e-09, 9.277076e-09, 9.273725e-09, 9.246322e-09, 9.274102e-09, 
    9.002945e-09, 8.995122e-09, 8.967964e-09, 8.989217e-09, 8.950494e-09, 
    8.972171e-09, 8.984634e-09, 9.032724e-09, 9.043289e-09, 9.053086e-09, 
    9.072435e-09, 9.097267e-09, 9.140829e-09, 9.178729e-09, 9.213328e-09, 
    9.210792e-09, 9.211685e-09, 9.219415e-09, 9.200269e-09, 9.222558e-09, 
    9.226299e-09, 9.216517e-09, 9.273276e-09, 9.257061e-09, 9.273654e-09, 
    9.263096e-09, 8.997665e-09, 9.010827e-09, 9.003715e-09, 9.017089e-09, 
    9.007668e-09, 9.049564e-09, 9.062125e-09, 9.120901e-09, 9.096778e-09, 
    9.135169e-09, 9.100678e-09, 9.10679e-09, 9.136423e-09, 9.102542e-09, 
    9.17664e-09, 9.126405e-09, 9.219715e-09, 9.169552e-09, 9.222858e-09, 
    9.213178e-09, 9.229205e-09, 9.24356e-09, 9.261618e-09, 9.294939e-09, 
    9.287223e-09, 9.315088e-09, 9.030448e-09, 9.047521e-09, 9.046017e-09, 
    9.063883e-09, 9.077096e-09, 9.105732e-09, 9.151662e-09, 9.13439e-09, 
    9.166097e-09, 9.172463e-09, 9.124292e-09, 9.153869e-09, 9.058946e-09, 
    9.074284e-09, 9.065151e-09, 9.031796e-09, 9.138371e-09, 9.083678e-09, 
    9.184672e-09, 9.155043e-09, 9.241513e-09, 9.19851e-09, 9.282975e-09, 
    9.319085e-09, 9.353066e-09, 9.392782e-09, 9.056838e-09, 9.045237e-09, 
    9.066008e-09, 9.094744e-09, 9.121405e-09, 9.15685e-09, 9.160477e-09, 
    9.167117e-09, 9.184316e-09, 9.198778e-09, 9.169217e-09, 9.202403e-09, 
    9.077842e-09, 9.143118e-09, 9.040853e-09, 9.071648e-09, 9.09305e-09, 
    9.083661e-09, 9.132416e-09, 9.143907e-09, 9.190603e-09, 9.166464e-09, 
    9.310174e-09, 9.246593e-09, 9.423018e-09, 9.373716e-09, 9.041185e-09, 
    9.056797e-09, 9.111135e-09, 9.085281e-09, 9.159216e-09, 9.177415e-09, 
    9.192209e-09, 9.211121e-09, 9.213162e-09, 9.224368e-09, 9.206006e-09, 
    9.223642e-09, 9.156926e-09, 9.186739e-09, 9.104923e-09, 9.124838e-09, 
    9.115676e-09, 9.105627e-09, 9.136641e-09, 9.169683e-09, 9.170388e-09, 
    9.180982e-09, 9.210841e-09, 9.159516e-09, 9.318383e-09, 9.220273e-09, 
    9.073822e-09, 9.103895e-09, 9.10819e-09, 9.09654e-09, 9.175591e-09, 
    9.146948e-09, 9.224094e-09, 9.203244e-09, 9.237406e-09, 9.220431e-09, 
    9.217933e-09, 9.19613e-09, 9.182556e-09, 9.148262e-09, 9.120358e-09, 
    9.09823e-09, 9.103375e-09, 9.127682e-09, 9.171704e-09, 9.213347e-09, 
    9.204226e-09, 9.23481e-09, 9.153855e-09, 9.187802e-09, 9.174682e-09, 
    9.208891e-09, 9.133932e-09, 9.197768e-09, 9.117614e-09, 9.124642e-09, 
    9.14638e-09, 9.190106e-09, 9.199777e-09, 9.210106e-09, 9.203732e-09, 
    9.172822e-09, 9.167756e-09, 9.145851e-09, 9.139804e-09, 9.123112e-09, 
    9.109294e-09, 9.121919e-09, 9.135179e-09, 9.172834e-09, 9.206768e-09, 
    9.243765e-09, 9.252818e-09, 9.296047e-09, 9.260859e-09, 9.318929e-09, 
    9.269561e-09, 9.355018e-09, 9.201465e-09, 9.268106e-09, 9.147368e-09, 
    9.160376e-09, 9.183903e-09, 9.237863e-09, 9.208731e-09, 9.242799e-09, 
    9.167557e-09, 9.128521e-09, 9.11842e-09, 9.099575e-09, 9.118851e-09, 
    9.117283e-09, 9.135727e-09, 9.1298e-09, 9.174084e-09, 9.150297e-09, 
    9.217871e-09, 9.24253e-09, 9.312169e-09, 9.354859e-09, 9.398313e-09, 
    9.417497e-09, 9.423337e-09, 9.425777e-09 ;

 H2OCAN =
  0.05992911, 0.05991415, 0.059917, 0.05990504, 0.05991156, 0.05990382, 
    0.05992595, 0.05991367, 0.05992144, 0.05992759, 0.05988215, 0.05990447, 
    0.05985781, 0.05987219, 0.05983553, 0.05986023, 0.05983046, 0.05983593, 
    0.05981864, 0.05982359, 0.05980198, 0.05981635, 0.05979019, 0.05980526, 
    0.05980302, 0.05981687, 0.05989969, 0.059885, 0.05990063, 0.05989852, 
    0.05989939, 0.05991154, 0.05991783, 0.05993005, 0.05992778, 0.05991869, 
    0.05989756, 0.05990455, 0.0598863, 0.0598867, 0.05986677, 0.05987577, 
    0.0598419, 0.0598515, 0.05982338, 0.05983053, 0.05982377, 0.05982578, 
    0.05982374, 0.05983421, 0.05982975, 0.05983883, 0.05987415, 0.0598639, 
    0.05989467, 0.05991368, 0.05992547, 0.05993403, 0.05993282, 0.05993058, 
    0.05991864, 0.0599071, 0.05989837, 0.05989255, 0.05988676, 0.05987026, 
    0.05986082, 0.05984011, 0.0598436, 0.05983747, 0.05983123, 0.05982107, 
    0.0598227, 0.05981828, 0.05983744, 0.05982482, 0.05984564, 0.05984, 
    0.05988625, 0.05990262, 0.05991044, 0.05991649, 0.05993192, 0.05992133, 
    0.05992553, 0.0599153, 0.05990892, 0.05991203, 0.05989239, 0.05990009, 
    0.05986026, 0.05987737, 0.05983195, 0.05984286, 0.05982929, 0.05983618, 
    0.05982446, 0.05983501, 0.05981654, 0.05981262, 0.05981532, 0.05980456, 
    0.05983562, 0.05982387, 0.05991217, 0.05991167, 0.05990921, 0.05992002, 
    0.05992062, 0.05993016, 0.05992157, 0.05991799, 0.05990847, 0.05990302, 
    0.05989775, 0.05988612, 0.05987346, 0.05985538, 0.05984217, 0.0598333, 
    0.05983867, 0.05983394, 0.05983927, 0.05984172, 0.05981416, 0.05982977, 
    0.05980612, 0.05980739, 0.05981821, 0.05980725, 0.0599113, 0.05991422, 
    0.05992464, 0.05991649, 0.05993118, 0.0599231, 0.05991852, 0.05990016, 
    0.05989585, 0.05989219, 0.0598847, 0.05987532, 0.05985888, 0.05984434, 
    0.05983082, 0.05983179, 0.05983146, 0.05982854, 0.05983591, 0.05982732, 
    0.05982597, 0.05982964, 0.05980757, 0.05981389, 0.05980742, 0.05981151, 
    0.05991324, 0.05990829, 0.05991098, 0.05990597, 0.05990959, 0.05989377, 
    0.05988901, 0.05986665, 0.05987556, 0.05986108, 0.05987401, 0.05987179, 
    0.05986105, 0.05987325, 0.05984534, 0.05986468, 0.05982842, 0.0598483, 
    0.0598272, 0.05983088, 0.05982467, 0.05981921, 0.05981213, 0.05979931, 
    0.05980224, 0.0597913, 0.05990079, 0.05989442, 0.05989479, 0.05988796, 
    0.05988301, 0.05987205, 0.05985465, 0.05986114, 0.059849, 0.05984662, 
    0.05986495, 0.0598539, 0.05989, 0.05988434, 0.05988755, 0.0599004, 
    0.05985991, 0.05988075, 0.05984198, 0.05985331, 0.05982002, 0.05983685, 
    0.0598039, 0.05979019, 0.05977627, 0.05976099, 0.05989072, 0.05989508, 
    0.0598871, 0.05987654, 0.05986617, 0.05985266, 0.05985117, 0.05984868, 
    0.059842, 0.05983645, 0.05984809, 0.05983504, 0.05988344, 0.05985801, 
    0.05989691, 0.05988539, 0.05987707, 0.05988052, 0.05986183, 0.05985748, 
    0.05983981, 0.05984885, 0.05979376, 0.05981834, 0.0597486, 0.05976844, 
    0.05989665, 0.05989064, 0.05987021, 0.05987987, 0.05985165, 0.05984475, 
    0.05983895, 0.05983184, 0.05983092, 0.05982666, 0.05983366, 0.05982687, 
    0.05985263, 0.05984113, 0.05987231, 0.05986486, 0.05986822, 0.05987205, 
    0.05986024, 0.05984795, 0.05984737, 0.05984348, 0.05983301, 0.05985153, 
    0.05979116, 0.05982921, 0.05988413, 0.05987313, 0.05987117, 0.05987551, 
    0.05984545, 0.05985642, 0.05982672, 0.05983472, 0.05982152, 0.05982812, 
    0.0598291, 0.05983747, 0.05984275, 0.05985598, 0.0598666, 0.05987484, 
    0.0598729, 0.05986383, 0.05984713, 0.05983098, 0.05983457, 0.05982252, 
    0.05985372, 0.05984086, 0.05984594, 0.0598326, 0.05986138, 0.05983786, 
    0.05986748, 0.05986482, 0.05985663, 0.0598402, 0.05983607, 0.05983223, 
    0.05983453, 0.05984664, 0.05984848, 0.05985675, 0.05985919, 0.05986538, 
    0.05987065, 0.05986591, 0.059861, 0.05984651, 0.05983354, 0.05981918, 
    0.05981553, 0.05979943, 0.05981299, 0.05979101, 0.05981038, 0.05977641, 
    0.05983602, 0.05981029, 0.05985615, 0.05985118, 0.05984251, 0.05982178, 
    0.05983266, 0.05981977, 0.05984852, 0.05986368, 0.0598672, 0.0598744, 
    0.05986703, 0.05986762, 0.05986057, 0.05986282, 0.05984602, 0.05985504, 
    0.05982921, 0.0598198, 0.05979257, 0.05977592, 0.05975832, 0.05975068, 
    0.05974832, 0.05974735 ;

 H2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO_TOP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSOI =
  3.844866, 3.857815, 3.855295, 3.86576, 3.859952, 3.866809, 3.847488, 
    3.85833, 3.851406, 3.84603, 3.886137, 3.866228, 3.906909, 3.894146, 
    3.926268, 3.904921, 3.930584, 3.925652, 3.940513, 3.93625, 3.955308, 
    3.942481, 3.965216, 3.952242, 3.954269, 3.942058, 3.870228, 3.883654, 
    3.869434, 3.871346, 3.870488, 3.860072, 3.854832, 3.843878, 3.845865, 
    3.853911, 3.872205, 3.865987, 3.881675, 3.88132, 3.898846, 3.890936, 
    3.920486, 3.912071, 3.936428, 3.930291, 3.93614, 3.934366, 3.936163, 
    3.927165, 3.931018, 3.923108, 3.892416, 3.901417, 3.874622, 3.858584, 
    3.847963, 3.840441, 3.841504, 3.84353, 3.853958, 3.863785, 3.871287, 
    3.876312, 3.881269, 3.896305, 3.904282, 3.922189, 3.918953, 3.924437, 
    3.929681, 3.938498, 3.937046, 3.940935, 3.924292, 3.935346, 3.917111, 
    3.922092, 3.882617, 3.867664, 3.861322, 3.855779, 3.842321, 3.851611, 
    3.847947, 3.856669, 3.86222, 3.859474, 3.87645, 3.869843, 3.904756, 
    3.889686, 3.929069, 3.919617, 3.931337, 3.925354, 3.935611, 3.926378, 
    3.942383, 3.945875, 3.943488, 3.952662, 3.925867, 3.93614, 3.859397, 
    3.859845, 3.861932, 3.852766, 3.852206, 3.843824, 3.851281, 3.854461, 
    3.862542, 3.867329, 3.871884, 3.881915, 3.893143, 3.908889, 3.92023, 
    3.927846, 3.923174, 3.927298, 3.922688, 3.920529, 3.944566, 3.931054, 
    3.951342, 3.950217, 3.941027, 3.950344, 3.860159, 3.857583, 3.848649, 
    3.855639, 3.842912, 3.850031, 3.85413, 3.86998, 3.873471, 3.876709, 
    3.883111, 3.89134, 3.905811, 3.918435, 3.929986, 3.929139, 3.929437, 
    3.932021, 3.925623, 3.933072, 3.934324, 3.931053, 3.950066, 3.944627, 
    3.950193, 3.946651, 3.85842, 3.862757, 3.860413, 3.864822, 3.861715, 
    3.875544, 3.879698, 3.899185, 3.891178, 3.903928, 3.892472, 3.8945, 
    3.904345, 3.89309, 3.917738, 3.901014, 3.932122, 3.915375, 3.933173, 
    3.929936, 3.935297, 3.940102, 3.946155, 3.957342, 3.954749, 3.96412, 
    3.86923, 3.874869, 3.874372, 3.88028, 3.884654, 3.894149, 3.909417, 
    3.90367, 3.914225, 3.916346, 3.900313, 3.910152, 3.878647, 3.883722, 
    3.8807, 3.869674, 3.904993, 3.886834, 3.920417, 3.910543, 3.939417, 
    3.925036, 3.953323, 3.965465, 3.97692, 3.99034, 3.877949, 3.874115, 
    3.880983, 3.890503, 3.899354, 3.911145, 3.912353, 3.914565, 3.920299, 
    3.925126, 3.915264, 3.926336, 3.8849, 3.906573, 3.872665, 3.88285, 
    3.889941, 3.886829, 3.903013, 3.906836, 3.922396, 3.914347, 3.962465, 
    3.941118, 4.000581, 3.983893, 3.872775, 3.877936, 3.895942, 3.887367, 
    3.911933, 3.917997, 3.922932, 3.929249, 3.929931, 3.933678, 3.92754, 
    3.933435, 3.91117, 3.921107, 3.893881, 3.900494, 3.897451, 3.894114, 
    3.904418, 3.915419, 3.915655, 3.919187, 3.929153, 3.912033, 3.965226, 
    3.932306, 3.88357, 3.893539, 3.894965, 3.891099, 3.917389, 3.907848, 
    3.933586, 3.926617, 3.938041, 3.932361, 3.931526, 3.924241, 3.919712, 
    3.908285, 3.899005, 3.89166, 3.893367, 3.901439, 3.916093, 3.929993, 
    3.926944, 3.937172, 3.910148, 3.921461, 3.917086, 3.928504, 3.903517, 
    3.924786, 3.898095, 3.900429, 3.907659, 3.92223, 3.925459, 3.92891, 
    3.92678, 3.916465, 3.914778, 3.907483, 3.90547, 3.899921, 3.895331, 
    3.899524, 3.903932, 3.91647, 3.927794, 3.940171, 3.943204, 3.957714, 
    3.945899, 3.96541, 3.948817, 3.977577, 3.926022, 3.94833, 3.907988, 
    3.912319, 3.92016, 3.938193, 3.92845, 3.939847, 3.914711, 3.901718, 
    3.898362, 3.892106, 3.898505, 3.897984, 3.904115, 3.902144, 3.916886, 
    3.908963, 3.931505, 3.939757, 3.963137, 3.977524, 3.992212, 3.99871, 
    4.00069, 4.001517,
  3.31989, 3.33258, 3.330112, 3.340366, 3.334677, 3.341394, 3.322462, 
    3.333082, 3.326301, 3.321034, 3.36033, 3.340825, 3.380714, 3.3682, 
    3.399711, 3.378761, 3.403949, 3.399112, 3.413702, 3.409518, 3.42822, 
    3.415635, 3.437957, 3.425215, 3.427203, 3.41522, 3.344749, 3.357895, 
    3.34397, 3.345842, 3.345003, 3.334792, 3.329651, 3.318926, 3.320872, 
    3.328753, 3.346684, 3.340593, 3.355974, 3.355626, 3.37281, 3.365054, 
    3.394042, 3.385786, 3.409693, 3.403667, 3.409408, 3.407667, 3.409431, 
    3.400598, 3.40438, 3.396617, 3.366504, 3.375331, 3.349055, 3.333325, 
    3.322926, 3.315558, 3.316599, 3.318583, 3.328799, 3.338434, 3.345789, 
    3.350715, 3.355576, 3.370306, 3.378137, 3.39571, 3.39254, 3.397917, 
    3.403068, 3.411723, 3.410298, 3.414114, 3.397779, 3.408627, 3.390733, 
    3.395619, 3.356877, 3.342236, 3.33601, 3.330585, 3.317399, 3.326499, 
    3.322909, 3.33146, 3.3369, 3.33421, 3.35085, 3.344372, 3.378602, 
    3.363824, 3.402467, 3.393191, 3.404694, 3.398822, 3.408887, 3.399827, 
    3.415537, 3.418963, 3.416621, 3.425632, 3.399325, 3.409406, 3.334133, 
    3.334572, 3.336618, 3.327631, 3.327083, 3.318871, 3.326179, 3.329293, 
    3.337217, 3.341908, 3.346373, 3.356207, 3.367214, 3.382659, 3.393791, 
    3.401268, 3.396683, 3.40073, 3.396205, 3.394087, 3.417678, 3.404414, 
    3.424335, 3.423231, 3.414204, 3.423355, 3.33488, 3.332356, 3.323599, 
    3.330451, 3.317979, 3.324952, 3.328966, 3.344502, 3.347929, 3.351102, 
    3.357381, 3.36545, 3.379641, 3.392028, 3.403369, 3.402537, 3.40283, 
    3.405365, 3.399085, 3.406397, 3.407623, 3.404415, 3.423083, 3.417741, 
    3.423207, 3.419729, 3.333177, 3.337426, 3.335129, 3.339449, 3.336404, 
    3.349955, 3.354027, 3.373138, 3.36529, 3.377793, 3.36656, 3.368547, 
    3.378192, 3.367168, 3.39134, 3.374929, 3.405463, 3.389016, 3.406496, 
    3.40332, 3.408582, 3.413297, 3.419241, 3.430224, 3.427679, 3.436883, 
    3.343771, 3.349296, 3.348814, 3.354605, 3.358893, 3.368206, 3.38318, 
    3.377544, 3.3879, 3.38998, 3.374252, 3.383899, 3.353001, 3.357974, 
    3.355015, 3.344205, 3.378836, 3.361026, 3.393975, 3.384285, 3.412624, 
    3.398504, 3.426278, 3.438195, 3.449459, 3.462636, 3.352319, 3.348561, 
    3.355296, 3.364624, 3.373309, 3.384875, 3.386063, 3.388232, 3.393861, 
    3.398597, 3.388914, 3.399786, 3.35912, 3.380388, 3.347137, 3.357117, 
    3.364075, 3.361026, 3.376902, 3.380651, 3.395914, 3.38802, 3.435247, 
    3.414289, 3.472709, 3.456303, 3.347248, 3.352308, 3.36996, 3.361553, 
    3.385651, 3.3916, 3.396446, 3.402642, 3.403314, 3.40699, 3.400967, 
    3.406754, 3.3849, 3.394653, 3.367944, 3.374427, 3.371445, 3.368173, 
    3.378279, 3.389065, 3.389302, 3.392765, 3.402527, 3.385749, 3.437947, 
    3.405625, 3.357832, 3.3676, 3.369005, 3.365216, 3.391003, 3.381641, 
    3.406902, 3.400062, 3.411276, 3.405699, 3.404879, 3.39773, 3.393283, 
    3.382069, 3.372967, 3.365766, 3.36744, 3.375353, 3.389727, 3.403372, 
    3.400378, 3.410423, 3.383899, 3.394998, 3.390702, 3.401912, 3.377393, 
    3.398244, 3.372077, 3.374366, 3.381456, 3.395747, 3.398925, 3.402309, 
    3.400222, 3.390094, 3.38844, 3.381285, 3.379308, 3.373868, 3.369366, 
    3.373477, 3.377798, 3.390101, 3.401213, 3.413364, 3.416345, 3.430578, 
    3.418979, 3.438127, 3.421829, 3.450087, 3.399465, 3.421364, 3.381781, 
    3.38603, 3.393718, 3.411417, 3.40186, 3.413042, 3.388376, 3.375623, 
    3.372338, 3.366202, 3.372479, 3.371968, 3.377981, 3.376049, 3.39051, 
    3.382737, 3.404857, 3.412955, 3.435915, 3.450046, 3.464486, 3.470873, 
    3.472819, 3.473632,
  3.010912, 3.024992, 3.022252, 3.033636, 3.027317, 3.034777, 3.013763, 
    3.025552, 3.018023, 3.012178, 3.055817, 3.034144, 3.078048, 3.064542, 
    3.098518, 3.075946, 3.103084, 3.097866, 3.113595, 3.109083, 3.129263, 
    3.115679, 3.139765, 3.126016, 3.128163, 3.115232, 3.038498, 3.053113, 
    3.037633, 3.039714, 3.03878, 3.027447, 3.021747, 3.009839, 3.011998, 
    3.020746, 3.04065, 3.033883, 3.050959, 3.050573, 3.069531, 3.061045, 
    3.092402, 3.083503, 3.109271, 3.102775, 3.108965, 3.107088, 3.10899, 
    3.099468, 3.103545, 3.095176, 3.062658, 3.072247, 3.04328, 3.025828, 
    3.014279, 3.006103, 3.007258, 3.00946, 3.020798, 3.031487, 3.03965, 
    3.04512, 3.050517, 3.066846, 3.075272, 3.094203, 3.090781, 3.09658, 
    3.10213, 3.111462, 3.109925, 3.114041, 3.096428, 3.108125, 3.088832, 
    3.0941, 3.051983, 3.035708, 3.028807, 3.022778, 3.008146, 3.018245, 
    3.014261, 3.023746, 3.029784, 3.026797, 3.04527, 3.038078, 3.075772, 
    3.059683, 3.101482, 3.091483, 3.103883, 3.097551, 3.108405, 3.098635, 
    3.115575, 3.119272, 3.116745, 3.126462, 3.098094, 3.108965, 3.026713, 
    3.0272, 3.02947, 3.019501, 3.018892, 3.009779, 3.017887, 3.021344, 
    3.030135, 3.035343, 3.0403, 3.05122, 3.063449, 3.080139, 3.09213, 
    3.100188, 3.095246, 3.099609, 3.094731, 3.092448, 3.117886, 3.103582, 
    3.125063, 3.123872, 3.114139, 3.124006, 3.027543, 3.02474, 3.015025, 
    3.022626, 3.008788, 3.016528, 3.020984, 3.038228, 3.042027, 3.045552, 
    3.052523, 3.061486, 3.076888, 3.090232, 3.102453, 3.101556, 3.101872, 
    3.104606, 3.097836, 3.105719, 3.107043, 3.103581, 3.123712, 3.117951, 
    3.123846, 3.120094, 3.025651, 3.030368, 3.027819, 3.032615, 3.029235, 
    3.044283, 3.048806, 3.069889, 3.061309, 3.074899, 3.062719, 3.064928, 
    3.075337, 3.063392, 3.089494, 3.07182, 3.104712, 3.086994, 3.105825, 
    3.1024, 3.108073, 3.11316, 3.119569, 3.13142, 3.128673, 3.138603, 
    3.037411, 3.043549, 3.043009, 3.04944, 3.054203, 3.064546, 3.080698, 
    3.074627, 3.08578, 3.088023, 3.071081, 3.081473, 3.047661, 3.053188, 
    3.049897, 3.037895, 3.076024, 3.056577, 3.092329, 3.081887, 3.112434, 
    3.097214, 3.127161, 3.140027, 3.152175, 3.166412, 3.046902, 3.042728, 
    3.050206, 3.060573, 3.070067, 3.082523, 3.0838, 3.086139, 3.092204, 
    3.09731, 3.086878, 3.098591, 3.05447, 3.077693, 3.04115, 3.052238, 
    3.059962, 3.056572, 3.073934, 3.077971, 3.094421, 3.085909, 3.136847, 
    3.114234, 3.177286, 3.159571, 3.04127, 3.046888, 3.066465, 3.057157, 
    3.083357, 3.089769, 3.09499, 3.101672, 3.102394, 3.106359, 3.099864, 
    3.106103, 3.08255, 3.093059, 3.064254, 3.071272, 3.068058, 3.064508, 
    3.075418, 3.087042, 3.087292, 3.091027, 3.101567, 3.083462, 3.139773, 
    3.104905, 3.053023, 3.06388, 3.065433, 3.061224, 3.089125, 3.07904, 
    3.106263, 3.098888, 3.110979, 3.104966, 3.104082, 3.096374, 3.091582, 
    3.079501, 3.0697, 3.061834, 3.063694, 3.07227, 3.087754, 3.102459, 
    3.099233, 3.110059, 3.08147, 3.093433, 3.088804, 3.100884, 3.074465, 
    3.096947, 3.068738, 3.071204, 3.07884, 3.094244, 3.097663, 3.101313, 
    3.09906, 3.088148, 3.086364, 3.078655, 3.076528, 3.070667, 3.065821, 
    3.070248, 3.074903, 3.088154, 3.100132, 3.113232, 3.116445, 3.131812, 
    3.119297, 3.139967, 3.122384, 3.152869, 3.098256, 3.121871, 3.079188, 
    3.083765, 3.092056, 3.111138, 3.100827, 3.112889, 3.086294, 3.072564, 
    3.069021, 3.06232, 3.069172, 3.068622, 3.075097, 3.073015, 3.088594, 
    3.080218, 3.104059, 3.112794, 3.137561, 3.152815, 3.168401, 3.1753, 
    3.177402, 3.178281,
  2.888639, 2.903944, 2.900963, 2.913344, 2.906471, 2.914585, 2.891737, 
    2.904553, 2.896366, 2.890014, 2.937405, 2.913897, 2.961275, 2.946599, 
    2.983575, 2.958987, 2.988553, 2.982863, 3.000012, 2.995091, 3.017113, 
    3.002285, 3.028578, 3.013566, 3.015911, 3.001797, 2.918632, 2.934543, 
    2.917691, 2.919955, 2.918939, 2.906613, 2.900417, 2.887471, 2.889818, 
    2.899328, 2.920974, 2.913611, 2.932193, 2.931772, 2.952, 2.942911, 
    2.976908, 2.967213, 2.995296, 2.988214, 2.994963, 2.992915, 2.99499, 
    2.984608, 2.989053, 2.97993, 2.944612, 2.954957, 2.923836, 2.904855, 
    2.892298, 2.883414, 2.884668, 2.887062, 2.899383, 2.911005, 2.919885, 
    2.925838, 2.931711, 2.949082, 2.958253, 2.978872, 2.975141, 2.981462, 
    2.98751, 2.997686, 2.996009, 3.0005, 2.981295, 2.994048, 2.973018, 
    2.978759, 2.933313, 2.915596, 2.908093, 2.901536, 2.885633, 2.896608, 
    2.892278, 2.902588, 2.909154, 2.905905, 2.926, 2.918175, 2.958797, 
    2.941476, 2.986804, 2.975907, 2.989421, 2.982518, 2.994353, 2.9837, 
    3.002172, 3.006207, 3.003449, 3.014052, 2.983111, 2.994963, 2.905814, 
    2.906343, 2.908812, 2.897974, 2.897311, 2.887407, 2.896218, 2.899977, 
    2.909534, 2.9152, 2.920593, 2.932477, 2.945448, 2.963551, 2.976612, 
    2.985393, 2.980006, 2.984761, 2.979446, 2.976957, 3.004695, 2.989094, 
    3.012525, 3.011225, 3.000607, 3.011371, 2.906715, 2.903668, 2.893108, 
    2.90137, 2.88633, 2.894742, 2.899587, 2.918339, 2.922471, 2.926307, 
    2.933895, 2.943376, 2.96001, 2.974545, 2.987862, 2.986885, 2.987229, 
    2.99021, 2.98283, 2.991423, 2.992867, 2.989092, 3.01105, 3.004764, 
    3.011197, 3.007102, 2.904658, 2.909789, 2.907016, 2.912232, 2.908556, 
    2.924928, 2.929851, 2.952392, 2.94319, 2.957845, 2.944676, 2.947006, 
    2.958325, 2.945386, 2.973742, 2.954495, 2.990326, 2.97102, 2.991539, 
    2.987804, 2.993989, 2.999538, 3.00653, 3.019465, 3.016466, 3.027308, 
    2.917449, 2.924128, 2.923539, 2.930539, 2.935699, 2.946602, 2.964159, 
    2.957547, 2.969694, 2.972137, 2.953686, 2.965004, 2.928604, 2.934621, 
    2.931037, 2.917976, 2.95907, 2.938203, 2.976828, 2.965454, 2.998747, 
    2.982153, 3.014816, 3.028867, 3.042136, 3.057704, 2.927777, 2.923234, 
    2.931373, 2.942415, 2.952584, 2.966147, 2.967537, 2.970085, 2.976692, 
    2.982256, 2.970891, 2.983652, 2.935984, 2.960887, 2.921518, 2.933587, 
    2.94177, 2.938196, 2.956792, 2.961189, 2.97911, 2.969834, 3.025394, 
    3.000712, 3.069598, 3.050222, 2.921648, 2.927761, 2.948663, 2.938812, 
    2.967054, 2.974039, 2.979727, 2.987011, 2.987798, 2.992122, 2.98504, 
    2.991842, 2.966176, 2.977623, 2.946294, 2.953895, 2.950396, 2.946562, 
    2.958408, 2.97107, 2.97134, 2.97541, 2.986905, 2.967169, 3.028594, 
    2.990542, 2.934439, 2.945903, 2.94754, 2.943099, 2.973339, 2.962353, 
    2.992016, 2.983976, 2.997159, 2.990602, 2.989638, 2.981236, 2.976015, 
    2.962856, 2.952184, 2.943743, 2.945704, 2.954982, 2.971846, 2.98787, 
    2.984354, 2.996155, 2.964999, 2.978032, 2.97299, 2.986152, 2.957371, 
    2.981868, 2.951136, 2.95382, 2.962135, 2.978918, 2.982641, 2.98662, 
    2.984164, 2.972275, 2.97033, 2.961933, 2.959618, 2.953236, 2.947961, 
    2.95278, 2.957849, 2.97228, 2.985333, 2.999617, 3.003121, 3.019897, 
    3.006236, 3.028807, 3.009611, 3.042901, 2.983291, 3.009046, 2.962514, 
    2.967499, 2.976533, 2.997335, 2.98609, 2.999244, 2.970254, 2.955303, 
    2.951444, 2.944255, 2.951608, 2.95101, 2.958058, 2.955791, 2.97276, 
    2.963635, 2.989614, 2.99914, 3.026171, 3.042837, 3.059876, 3.067423, 
    3.069723, 3.070685,
  2.94331, 2.959417, 2.956279, 2.969319, 2.962078, 2.970627, 2.946568, 
    2.960059, 2.951439, 2.944756, 2.994787, 2.969902, 3.020844, 3.004816, 
    3.045234, 3.018345, 3.050683, 3.044453, 3.063145, 3.057845, 3.081308, 
    3.065558, 3.093498, 3.077538, 3.08003, 3.06504, 2.974892, 2.991678, 
    2.973901, 2.976288, 2.975216, 2.962228, 2.955704, 2.942082, 2.94455, 
    2.954557, 2.977362, 2.969601, 2.989196, 2.988752, 3.010713, 3.000792, 
    3.037936, 3.027333, 3.05807, 3.050312, 3.057706, 3.055462, 3.057735, 
    3.046364, 3.051231, 3.041244, 3.002648, 3.013942, 2.98038, 2.960377, 
    2.947159, 2.937815, 2.939134, 2.941651, 2.954616, 2.966854, 2.976214, 
    2.982491, 2.988688, 3.007527, 3.017542, 3.040086, 3.036004, 3.042921, 
    3.049541, 3.060678, 3.058852, 3.063663, 3.042737, 3.056703, 3.033681, 
    3.039961, 2.990381, 2.971693, 2.963788, 2.956882, 2.940149, 2.951695, 
    2.947138, 2.957989, 2.964904, 2.961482, 2.982663, 2.974411, 3.018137, 
    2.999226, 3.048768, 3.036841, 3.051634, 3.044076, 3.057037, 3.04537, 
    3.065438, 3.069721, 3.066794, 3.078054, 3.044725, 3.057706, 2.961386, 
    2.961944, 2.964544, 2.953132, 2.952435, 2.942014, 2.951284, 2.95524, 
    2.965305, 2.971275, 2.97696, 2.989497, 3.00356, 3.023331, 3.037613, 
    3.047223, 3.041326, 3.046532, 3.040714, 3.03799, 3.068116, 3.051277, 
    3.076432, 3.07505, 3.063777, 3.075206, 2.962336, 2.959126, 2.948011, 
    2.956706, 2.940881, 2.94973, 2.95483, 2.974584, 2.97894, 2.982987, 
    2.990993, 3.001299, 3.019462, 3.035351, 3.049927, 3.048856, 3.049233, 
    3.052498, 3.044417, 3.053827, 3.055409, 3.051274, 3.074865, 3.068189, 
    3.075021, 3.070672, 2.960169, 2.965573, 2.962652, 2.968148, 2.964275, 
    2.981533, 2.986726, 3.011141, 3.001096, 3.017096, 3.002717, 3.00526, 
    3.017622, 3.003492, 3.034474, 3.013438, 3.052625, 3.031498, 3.053954, 
    3.049863, 3.056639, 3.062643, 3.070064, 3.083807, 3.080619, 3.092148, 
    2.973646, 2.980688, 2.980067, 2.987452, 2.992925, 3.00482, 3.023995, 
    3.01677, 3.030046, 3.032718, 3.012553, 3.02492, 2.98541, 2.99176, 
    2.987977, 2.974202, 3.018435, 2.995656, 3.03785, 3.025411, 3.061803, 
    3.043677, 3.078866, 3.093806, 3.10793, 3.124524, 2.984538, 2.979745, 
    2.988331, 3.000251, 3.01135, 3.026168, 3.027688, 3.030474, 3.0377, 
    3.043789, 3.031356, 3.045317, 2.993237, 3.02042, 2.977936, 2.990669, 
    2.999547, 2.995648, 3.015945, 3.020749, 3.040346, 3.030199, 3.090113, 
    3.063889, 3.137215, 3.116547, 2.978072, 2.98452, 3.00707, 2.99632, 
    3.02716, 3.034798, 3.041021, 3.048995, 3.049857, 3.054592, 3.046836, 
    3.054285, 3.0262, 3.038719, 3.004483, 3.012782, 3.008961, 3.004776, 
    3.01771, 3.031552, 3.031846, 3.036299, 3.048881, 3.027285, 3.093517, 
    3.052865, 2.991567, 3.004057, 3.005843, 3.000996, 3.034032, 3.022021, 
    3.054477, 3.045671, 3.060111, 3.052928, 3.051872, 3.042673, 3.03696, 
    3.022571, 3.010913, 3.001698, 3.003839, 3.013969, 3.0324, 3.049936, 
    3.046086, 3.059011, 3.024913, 3.039167, 3.033651, 3.048054, 3.016579, 
    3.043367, 3.009769, 3.0127, 3.021783, 3.040137, 3.04421, 3.048567, 
    3.045877, 3.032869, 3.030742, 3.021562, 3.019033, 3.012061, 3.006302, 
    3.011564, 3.0171, 3.032874, 3.047158, 3.062726, 3.066445, 3.084268, 
    3.069753, 3.093744, 3.073339, 3.108747, 3.044924, 3.072738, 3.022197, 
    3.027646, 3.037527, 3.060306, 3.047986, 3.062331, 3.030659, 3.01432, 
    3.010104, 3.002258, 3.010284, 3.00963, 3.017328, 3.014853, 3.033399, 
    3.023423, 3.051846, 3.062221, 3.090938, 3.108678, 3.12684, 3.134893, 
    3.137349, 3.138376,
  2.96992, 2.988319, 2.984731, 2.999652, 2.991363, 3.00115, 2.973638, 
    2.989053, 2.979201, 2.971569, 3.028873, 3.000319, 3.058882, 3.04041, 
    3.087076, 3.055999, 3.09339, 3.086172, 3.107955, 3.101695, 3.129773, 
    3.11085, 3.144451, 3.125239, 3.128236, 3.110228, 3.006037, 3.025301, 
    3.004901, 3.007638, 3.006409, 2.991534, 2.984074, 2.968518, 2.971334, 
    2.982763, 3.008869, 2.999974, 3.022449, 3.021939, 3.047201, 3.035779, 
    3.078629, 3.066374, 3.101956, 3.092959, 3.101533, 3.098929, 3.101567, 
    3.088385, 3.094024, 3.082456, 3.037914, 3.050922, 3.01233, 2.989418, 
    2.974312, 2.963651, 2.965156, 2.968026, 2.98283, 2.996829, 3.007552, 
    3.014751, 3.021866, 3.043532, 3.055073, 3.081116, 3.076394, 3.084398, 
    3.092066, 3.104996, 3.102863, 3.108577, 3.084185, 3.100369, 3.073709, 
    3.080972, 3.02381, 3.002371, 2.99332, 2.98542, 2.966313, 2.979493, 
    2.974289, 2.986686, 2.994597, 2.990681, 3.014949, 3.005486, 3.055759, 
    3.033978, 3.09117, 3.077362, 3.094491, 3.085735, 3.100757, 3.087234, 
    3.110706, 3.115848, 3.112333, 3.125859, 3.086486, 3.101533, 2.990571, 
    2.99121, 2.994185, 2.981134, 2.980338, 2.968441, 2.979023, 2.983544, 
    2.995056, 3.001892, 3.008407, 3.022794, 3.038964, 3.061753, 3.078255, 
    3.08938, 3.082552, 3.088579, 3.081843, 3.078691, 3.11392, 3.094077, 
    3.123909, 3.122248, 3.108713, 3.122436, 2.991658, 2.987987, 2.975285, 
    2.98522, 2.967149, 2.977248, 2.983075, 3.005684, 3.010679, 3.015321, 
    3.024513, 3.036362, 3.057287, 3.075639, 3.092512, 3.091272, 3.091708, 
    3.095493, 3.08613, 3.097034, 3.098869, 3.094074, 3.122026, 3.114008, 
    3.122213, 3.116989, 2.989179, 2.995363, 2.99202, 2.99831, 2.993877, 
    3.013652, 3.019612, 3.047694, 3.036129, 3.054559, 3.037994, 3.040921, 
    3.055165, 3.038886, 3.074625, 3.050341, 3.09564, 3.071185, 3.097181, 
    3.092439, 3.100295, 3.107352, 3.116259, 3.13278, 3.128944, 3.142823, 
    3.004609, 3.012683, 3.01197, 3.020446, 3.026733, 3.040414, 3.062519, 
    3.054183, 3.069507, 3.072595, 3.049322, 3.063586, 3.018101, 3.025394, 
    3.021049, 3.005246, 3.056103, 3.029872, 3.078529, 3.064153, 3.106345, 
    3.085273, 3.126835, 3.144822, 3.161329, 3.180762, 3.0171, 3.011601, 
    3.021455, 3.035156, 3.047935, 3.065028, 3.066783, 3.070001, 3.078356, 
    3.085402, 3.071021, 3.087172, 3.027092, 3.058392, 3.009526, 3.02414, 
    3.034346, 3.029863, 3.053231, 3.058772, 3.081417, 3.069684, 3.140372, 
    3.108848, 3.195661, 3.171414, 3.009683, 3.017081, 3.043005, 3.030636, 
    3.066173, 3.075, 3.082199, 3.091433, 3.092432, 3.097921, 3.088932, 
    3.097565, 3.065065, 3.079535, 3.040026, 3.049585, 3.045182, 3.040363, 
    3.055267, 3.071247, 3.071588, 3.076735, 3.091301, 3.066318, 3.144474, 
    3.095918, 3.025173, 3.039536, 3.041592, 3.036014, 3.074114, 3.060241, 
    3.097787, 3.087583, 3.104324, 3.095991, 3.094767, 3.08411, 3.0775, 
    3.060876, 3.047431, 3.036822, 3.039284, 3.050953, 3.072228, 3.092523, 
    3.088063, 3.103048, 3.063579, 3.080053, 3.073673, 3.090343, 3.053962, 
    3.084914, 3.046113, 3.04949, 3.059966, 3.081176, 3.08589, 3.090937, 
    3.087821, 3.07277, 3.070312, 3.059711, 3.056792, 3.048754, 3.04212, 
    3.048182, 3.054563, 3.072775, 3.089305, 3.107453, 3.111914, 3.133334, 
    3.115886, 3.144748, 3.120193, 3.162284, 3.086717, 3.11947, 3.060443, 
    3.066734, 3.078156, 3.104551, 3.090264, 3.106979, 3.070215, 3.051358, 
    3.0465, 3.037466, 3.046707, 3.045954, 3.054826, 3.051972, 3.073382, 
    3.061858, 3.094737, 3.106846, 3.141365, 3.162204, 3.183479, 3.192933, 
    3.195818, 3.197025,
  3.254737, 3.278214, 3.273626, 3.292734, 3.282109, 3.294657, 3.259472, 
    3.279153, 3.266564, 3.256837, 3.3299, 3.29359, 3.367675, 3.344384, 
    3.40347, 3.364032, 3.411527, 3.402317, 3.430173, 3.422149, 3.458259, 
    3.433888, 3.477261, 3.452407, 3.456274, 3.43309, 3.300935, 3.325425, 
    3.299475, 3.302993, 3.301413, 3.282329, 3.272787, 3.252954, 3.256538, 
    3.271112, 3.304577, 3.293148, 3.321856, 3.321218, 3.352931, 3.338563, 
    3.392715, 3.377157, 3.422483, 3.410977, 3.421941, 3.418609, 3.421985, 
    3.405139, 3.412338, 3.397584, 3.341246, 3.357622, 3.309032, 3.279619, 
    3.260331, 3.246767, 3.248678, 3.252328, 3.271198, 3.289113, 3.302883, 
    3.312152, 3.321126, 3.348311, 3.362862, 3.395878, 3.389873, 3.400056, 
    3.409836, 3.426378, 3.423645, 3.43097, 3.399785, 3.420452, 3.386461, 
    3.395695, 3.323559, 3.296224, 3.284615, 3.274507, 3.250149, 3.266937, 
    3.260301, 3.276125, 3.286251, 3.281236, 3.312406, 3.300226, 3.363728, 
    3.336303, 3.408693, 3.391104, 3.412934, 3.401761, 3.420948, 3.403671, 
    3.433704, 3.440311, 3.435794, 3.453207, 3.402718, 3.421942, 3.281096, 
    3.281913, 3.285723, 3.269032, 3.268015, 3.252856, 3.266338, 3.27211, 
    3.286839, 3.295609, 3.303983, 3.322288, 3.342566, 3.371306, 3.392239, 
    3.406408, 3.397706, 3.405386, 3.396803, 3.392793, 3.437833, 3.412405, 
    3.450692, 3.448552, 3.431145, 3.448793, 3.282487, 3.277789, 3.261571, 
    3.274251, 3.251212, 3.264074, 3.27151, 3.300481, 3.306906, 3.312885, 
    3.324439, 3.339296, 3.365659, 3.388914, 3.410406, 3.408823, 3.40938, 
    3.414215, 3.402264, 3.416184, 3.418532, 3.412401, 3.448265, 3.437946, 
    3.448506, 3.44178, 3.279314, 3.287233, 3.28295, 3.291012, 3.285329, 
    3.310735, 3.318309, 3.353553, 3.339003, 3.362213, 3.341346, 3.345027, 
    3.362978, 3.342467, 3.387626, 3.35689, 3.414403, 3.383258, 3.416373, 
    3.410313, 3.420356, 3.4294, 3.44084, 3.462145, 3.457189, 3.475149, 
    3.299099, 3.309487, 3.308569, 3.31935, 3.327218, 3.344388, 3.372275, 
    3.361737, 3.381129, 3.385048, 3.355605, 3.373627, 3.31642, 3.325542, 
    3.320105, 3.299917, 3.364163, 3.331152, 3.392587, 3.374345, 3.428108, 
    3.401172, 3.454467, 3.477742, 3.499918, 3.526191, 3.31517, 3.308093, 
    3.320613, 3.337782, 3.353856, 3.375453, 3.377676, 3.381756, 3.392366, 
    3.401337, 3.38305, 3.403592, 3.327668, 3.367056, 3.305423, 3.323972, 
    3.336765, 3.331141, 3.360537, 3.367536, 3.396261, 3.381354, 3.471971, 
    3.431318, 3.546055, 3.513531, 3.305624, 3.315145, 3.347648, 3.33211, 
    3.376903, 3.388102, 3.397256, 3.409029, 3.410303, 3.41732, 3.405836, 
    3.416864, 3.375499, 3.393867, 3.343901, 3.355936, 3.350389, 3.344325, 
    3.363107, 3.383337, 3.383769, 3.390306, 3.408861, 3.377086, 3.477291, 
    3.414758, 3.325265, 3.343285, 3.34587, 3.338859, 3.386976, 3.369393, 
    3.417148, 3.404116, 3.425517, 3.414851, 3.413287, 3.399691, 3.391278, 
    3.370196, 3.353222, 3.339874, 3.342969, 3.357662, 3.384581, 3.41042, 
    3.404728, 3.423882, 3.373617, 3.394526, 3.386416, 3.407636, 3.361459, 
    3.400715, 3.351561, 3.355817, 3.369046, 3.395954, 3.401958, 3.408395, 
    3.40442, 3.385269, 3.38215, 3.368722, 3.365034, 3.35489, 3.346535, 
    3.354167, 3.362218, 3.385276, 3.406312, 3.429529, 3.435256, 3.462861, 
    3.440361, 3.477646, 3.445904, 3.501205, 3.403012, 3.444973, 3.369649, 
    3.377614, 3.392113, 3.425807, 3.407536, 3.428921, 3.382028, 3.358173, 
    3.352048, 3.340683, 3.352309, 3.351361, 3.36255, 3.358947, 3.386047, 
    3.371439, 3.413249, 3.428751, 3.473259, 3.501097, 3.529877, 3.542453, 
    3.546262, 3.547857,
  3.812393, 3.852924, 3.844952, 3.878324, 3.859713, 3.881707, 3.820515, 
    3.854559, 3.83273, 3.815992, 3.945428, 3.879831, 4.016906, 3.972589, 
    4.084889, 4.009922, 4.10039, 4.08268, 4.136661, 4.120983, 4.192374, 
    4.143956, 4.230834, 4.180657, 4.188393, 4.142387, 3.892786, 3.937095, 
    3.890204, 3.896427, 3.893631, 3.860096, 3.843496, 3.80934, 3.815479, 
    3.840593, 3.899234, 3.879051, 3.93047, 3.929288, 3.98876, 3.961638, 
    4.064354, 4.034962, 4.121634, 4.099329, 4.120579, 4.114101, 4.120664, 
    4.088092, 4.101956, 4.073629, 3.96668, 3.997681, 3.907147, 3.855371, 
    3.821991, 3.798779, 3.802037, 3.808271, 3.840742, 3.871965, 3.896233, 
    3.912702, 3.929118, 3.980006, 4.007683, 4.070376, 4.058958, 4.078352, 
    4.097129, 4.129234, 4.123899, 4.138225, 4.077834, 4.117682, 4.052496, 
    4.070027, 3.933629, 3.884468, 3.86409, 3.846481, 3.804548, 3.833373, 
    3.82194, 3.849291, 3.866952, 3.858189, 3.913155, 3.891532, 4.00934, 
    3.957397, 4.094926, 4.061294, 4.103108, 4.081614, 4.118647, 4.085274, 
    4.143593, 4.15662, 4.147705, 4.182254, 4.083447, 4.120581, 3.857945, 
    3.85937, 3.866028, 3.836994, 3.835236, 3.809173, 3.832339, 3.842322, 
    3.867982, 3.883384, 3.898182, 3.931272, 3.969163, 4.023888, 4.063449, 
    4.09053, 4.073862, 4.088567, 4.072139, 4.064504, 4.151726, 4.102087, 
    4.177233, 4.172968, 4.138568, 4.173448, 3.860372, 3.852184, 3.824124, 
    3.846035, 3.806363, 3.828434, 3.841284, 3.891984, 3.903367, 3.91401, 
    3.935263, 3.963014, 4.01304, 4.05714, 4.098228, 4.095176, 4.09625, 
    4.105584, 4.082578, 4.109397, 4.113951, 4.102079, 4.172398, 4.151948, 
    4.172877, 4.159524, 3.85484, 3.86867, 3.86118, 3.875299, 3.865338, 
    3.910178, 3.923903, 3.98994, 3.962463, 4.006441, 3.966868, 3.973802, 
    4.007905, 3.968978, 4.054699, 3.996286, 4.105948, 4.046445, 4.109763, 
    4.098048, 4.117496, 4.135146, 4.157666, 4.200188, 4.190227, 4.226528, 
    3.889541, 3.907957, 3.906323, 3.925829, 3.940431, 3.972598, 4.025756, 
    4.005533, 4.042431, 4.049824, 3.99384, 4.028343, 3.920414, 3.937313, 
    3.927225, 3.890987, 4.010172, 3.947763, 4.064112, 4.029688, 4.132616, 
    4.080487, 4.184773, 4.231818, 4.277537, 4.332245, 3.918106, 3.905478, 
    3.928166, 3.960172, 3.990517, 4.031764, 4.035936, 4.043613, 4.063693, 
    4.080802, 4.046052, 4.085124, 3.941267, 4.015718, 3.900735, 3.934397, 
    3.958264, 3.947742, 4.003239, 4.01664, 4.071106, 4.042855, 4.220065, 
    4.138907, 4.374605, 4.306057, 3.901093, 3.918061, 3.978752, 3.949552, 
    4.034484, 4.055602, 4.073004, 4.095573, 4.09803, 4.111598, 4.089432, 
    4.110715, 4.031851, 4.066545, 3.971678, 3.994471, 3.983939, 3.972478, 
    4.008152, 4.046594, 4.047409, 4.05978, 4.095249, 4.034829, 4.230896, 
    4.106637, 3.936798, 3.970517, 3.975393, 3.962193, 4.05347, 4.020208, 
    4.111265, 4.086128, 4.127552, 4.106816, 4.103791, 4.077653, 4.061625, 
    4.021752, 3.989313, 3.964099, 3.969922, 3.997757, 4.048942, 4.098255, 
    4.087304, 4.124361, 4.028325, 4.067799, 4.052412, 4.092893, 4.005001, 
    4.079612, 3.986161, 3.994244, 4.01954, 4.070521, 4.081992, 4.094354, 
    4.086711, 4.050242, 4.044355, 4.018919, 4.011841, 3.99248, 3.976649, 
    3.991108, 4.006452, 4.050255, 4.090346, 4.1354, 4.146646, 4.201631, 
    4.156718, 4.231621, 4.167703, 4.280221, 4.084011, 4.165854, 4.0207, 
    4.03582, 4.06321, 4.128119, 4.0927, 4.134209, 4.044124, 3.998729, 
    3.987085, 3.96562, 3.98758, 3.985781, 4.007087, 4.000206, 4.051712, 
    4.024145, 4.103716, 4.133875, 4.222682, 4.279995, 4.339895, 4.366773, 
    4.375056, 4.378533,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HC =
  24814.08, 24834.51, 24830.5, 24847.23, 24837.91, 24848.92, 24818.18, 
    24835.33, 24824.35, 24815.9, 24880.44, 24847.98, 24915.19, 24893.71, 
    24948.14, 24911.82, 24955.61, 24947.08, 24972.99, 24965.5, 24999.43, 
    24976.47, 25017.51, 24993.89, 24997.54, 24975.72, 24854.44, 24876.36, 
    24853.16, 24856.26, 24854.86, 24838.11, 24829.77, 24812.53, 24815.64, 
    24828.31, 24857.65, 24847.59, 24873.11, 24872.52, 24901.57, 24888.37, 
    24938.22, 24923.94, 24965.81, 24955.1, 24965.3, 24962.2, 24965.35, 
    24949.69, 24956.37, 24942.71, 24890.83, 24905.89, 24861.59, 24835.74, 
    24818.93, 24807.18, 24808.83, 24811.99, 24828.38, 24844.05, 24856.16, 
    24864.34, 24872.44, 24897.32, 24910.74, 24941.13, 24935.6, 24944.99, 
    24954.04, 24969.45, 24966.89, 24973.74, 24944.74, 24963.92, 24932.47, 
    24940.96, 24874.66, 24850.29, 24840.11, 24831.27, 24810.1, 24824.67, 
    24818.9, 24832.68, 24841.54, 24837.15, 24864.57, 24853.82, 24911.54, 
    24886.3, 24952.98, 24936.73, 24956.92, 24946.56, 24964.38, 24948.33, 
    24976.3, 24982.49, 24978.25, 24994.64, 24947.45, 24965.3, 24837.03, 
    24837.74, 24841.08, 24826.5, 24825.61, 24812.45, 24824.15, 24829.18, 
    24842.06, 24849.75, 24857.13, 24873.5, 24892.04, 24918.56, 24937.78, 
    24950.87, 24942.82, 24949.92, 24941.99, 24938.29, 24980.17, 24956.43, 
    24992.27, 24990.25, 24973.9, 24990.48, 24838.24, 24834.14, 24820.01, 
    24831.05, 24811.02, 24822.18, 24828.66, 24854.04, 24859.71, 24864.99, 
    24875.46, 24889.04, 24913.33, 24934.72, 24954.57, 24953.1, 24953.62, 
    24958.11, 24947.03, 24959.94, 24962.13, 24956.42, 24989.98, 24980.27, 
    24990.21, 24983.87, 24835.47, 24842.4, 24838.65, 24845.72, 24840.73, 
    24863.09, 24869.88, 24902.14, 24888.77, 24910.14, 24890.92, 24894.3, 
    24910.84, 24891.95, 24933.54, 24905.22, 24958.29, 24929.53, 24960.12, 
    24954.49, 24963.83, 24972.27, 24982.99, 25003.11, 24998.41, 25015.49, 
    24852.83, 24861.99, 24861.18, 24870.82, 24878, 24893.71, 24919.46, 
    24909.7, 24927.58, 24931.17, 24904.03, 24920.71, 24868.16, 24876.47, 
    24871.51, 24853.55, 24911.94, 24881.59, 24938.1, 24921.37, 24971.06, 
    24946.02, 24995.84, 25017.97, 25039.25, 25064.59, 24867.02, 24860.76, 
    24871.97, 24887.65, 24902.42, 24922.38, 24924.41, 24928.15, 24937.9, 
    24946.17, 24929.34, 24948.26, 24878.4, 24914.62, 24858.4, 24875.04, 
    24886.72, 24881.58, 24908.59, 24915.06, 24941.49, 24927.78, 25012.46, 
    24974.06, 25084.1, 25052.43, 24858.58, 24867, 24896.71, 24882.46, 
    24923.71, 24933.97, 24942.4, 24953.29, 24954.48, 24961, 24950.34, 
    24960.57, 24922.42, 24939.28, 24893.26, 24904.34, 24899.23, 24893.65, 
    24910.96, 24929.6, 24930, 24936, 24953.14, 24923.88, 25017.54, 24958.62, 
    24876.21, 24892.7, 24895.07, 24888.64, 24932.94, 24916.79, 24960.84, 
    24948.74, 24968.64, 24958.7, 24957.25, 24944.65, 24936.9, 24917.53, 
    24901.84, 24889.57, 24892.41, 24905.93, 24930.74, 24954.58, 24949.31, 
    24967.12, 24920.7, 24939.89, 24932.43, 24952, 24909.44, 24945.6, 
    24900.31, 24904.23, 24916.46, 24941.2, 24946.75, 24952.71, 24949.02, 
    24931.37, 24928.51, 24916.16, 24912.75, 24903.37, 24895.68, 24902.71, 
    24910.14, 24931.38, 24950.78, 24972.39, 24977.75, 25003.79, 24982.54, 
    25017.88, 24987.75, 25040.49, 24947.72, 24986.88, 24917.03, 24924.36, 
    24937.66, 24968.91, 24951.91, 24971.82, 24928.4, 24906.4, 24900.76, 
    24890.31, 24901, 24900.12, 24910.45, 24907.12, 24932.09, 24918.69, 
    24957.21, 24971.66, 25013.69, 25040.38, 25068.13, 25080.51, 25084.3, 
    25085.9 ;

 HCSOI =
  24814.08, 24834.51, 24830.5, 24847.23, 24837.91, 24848.92, 24818.18, 
    24835.33, 24824.35, 24815.9, 24880.44, 24847.98, 24915.19, 24893.71, 
    24948.14, 24911.82, 24955.61, 24947.08, 24972.99, 24965.5, 24999.43, 
    24976.47, 25017.51, 24993.89, 24997.54, 24975.72, 24854.44, 24876.36, 
    24853.16, 24856.26, 24854.86, 24838.11, 24829.77, 24812.53, 24815.64, 
    24828.31, 24857.65, 24847.59, 24873.11, 24872.52, 24901.57, 24888.37, 
    24938.22, 24923.94, 24965.81, 24955.1, 24965.3, 24962.2, 24965.35, 
    24949.69, 24956.37, 24942.71, 24890.83, 24905.89, 24861.59, 24835.74, 
    24818.93, 24807.18, 24808.83, 24811.99, 24828.38, 24844.05, 24856.16, 
    24864.34, 24872.44, 24897.32, 24910.74, 24941.13, 24935.6, 24944.99, 
    24954.04, 24969.45, 24966.89, 24973.74, 24944.74, 24963.92, 24932.47, 
    24940.96, 24874.66, 24850.29, 24840.11, 24831.27, 24810.1, 24824.67, 
    24818.9, 24832.68, 24841.54, 24837.15, 24864.57, 24853.82, 24911.54, 
    24886.3, 24952.98, 24936.73, 24956.92, 24946.56, 24964.38, 24948.33, 
    24976.3, 24982.49, 24978.25, 24994.64, 24947.45, 24965.3, 24837.03, 
    24837.74, 24841.08, 24826.5, 24825.61, 24812.45, 24824.15, 24829.18, 
    24842.06, 24849.75, 24857.13, 24873.5, 24892.04, 24918.56, 24937.78, 
    24950.87, 24942.82, 24949.92, 24941.99, 24938.29, 24980.17, 24956.43, 
    24992.27, 24990.25, 24973.9, 24990.48, 24838.24, 24834.14, 24820.01, 
    24831.05, 24811.02, 24822.18, 24828.66, 24854.04, 24859.71, 24864.99, 
    24875.46, 24889.04, 24913.33, 24934.72, 24954.57, 24953.1, 24953.62, 
    24958.11, 24947.03, 24959.94, 24962.13, 24956.42, 24989.98, 24980.27, 
    24990.21, 24983.87, 24835.47, 24842.4, 24838.65, 24845.72, 24840.73, 
    24863.09, 24869.88, 24902.14, 24888.77, 24910.14, 24890.92, 24894.3, 
    24910.84, 24891.95, 24933.54, 24905.22, 24958.29, 24929.53, 24960.12, 
    24954.49, 24963.83, 24972.27, 24982.99, 25003.11, 24998.41, 25015.49, 
    24852.83, 24861.99, 24861.18, 24870.82, 24878, 24893.71, 24919.46, 
    24909.7, 24927.58, 24931.17, 24904.03, 24920.71, 24868.16, 24876.47, 
    24871.51, 24853.55, 24911.94, 24881.59, 24938.1, 24921.37, 24971.06, 
    24946.02, 24995.84, 25017.97, 25039.25, 25064.59, 24867.02, 24860.76, 
    24871.97, 24887.65, 24902.42, 24922.38, 24924.41, 24928.15, 24937.9, 
    24946.17, 24929.34, 24948.26, 24878.4, 24914.62, 24858.4, 24875.04, 
    24886.72, 24881.58, 24908.59, 24915.06, 24941.49, 24927.78, 25012.46, 
    24974.06, 25084.1, 25052.43, 24858.58, 24867, 24896.71, 24882.46, 
    24923.71, 24933.97, 24942.4, 24953.29, 24954.48, 24961, 24950.34, 
    24960.57, 24922.42, 24939.28, 24893.26, 24904.34, 24899.23, 24893.65, 
    24910.96, 24929.6, 24930, 24936, 24953.14, 24923.88, 25017.54, 24958.62, 
    24876.21, 24892.7, 24895.07, 24888.64, 24932.94, 24916.79, 24960.84, 
    24948.74, 24968.64, 24958.7, 24957.25, 24944.65, 24936.9, 24917.53, 
    24901.84, 24889.57, 24892.41, 24905.93, 24930.74, 24954.58, 24949.31, 
    24967.12, 24920.7, 24939.89, 24932.43, 24952, 24909.44, 24945.6, 
    24900.31, 24904.23, 24916.46, 24941.2, 24946.75, 24952.71, 24949.02, 
    24931.37, 24928.51, 24916.16, 24912.75, 24903.37, 24895.68, 24902.71, 
    24910.14, 24931.38, 24950.78, 24972.39, 24977.75, 25003.79, 24982.54, 
    25017.88, 24987.75, 25040.49, 24947.72, 24986.88, 24917.03, 24924.36, 
    24937.66, 24968.91, 24951.91, 24971.82, 24928.4, 24906.4, 24900.76, 
    24890.31, 24901, 24900.12, 24910.45, 24907.12, 24932.09, 24918.69, 
    24957.21, 24971.66, 25013.69, 25040.38, 25068.13, 25080.51, 25084.3, 
    25085.9 ;

 HEAT_FROM_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HR =
  6.35757e-08, 6.385525e-08, 6.38009e-08, 6.402639e-08, 6.39013e-08, 
    6.404895e-08, 6.363237e-08, 6.386636e-08, 6.371699e-08, 6.360087e-08, 
    6.446398e-08, 6.403645e-08, 6.490803e-08, 6.463537e-08, 6.532027e-08, 
    6.48656e-08, 6.541195e-08, 6.530715e-08, 6.562256e-08, 6.55322e-08, 
    6.593564e-08, 6.566426e-08, 6.614476e-08, 6.587083e-08, 6.591368e-08, 
    6.565531e-08, 6.412248e-08, 6.441076e-08, 6.41054e-08, 6.41465e-08, 
    6.412806e-08, 6.390389e-08, 6.379094e-08, 6.355432e-08, 6.359728e-08, 
    6.377105e-08, 6.416499e-08, 6.403126e-08, 6.436827e-08, 6.436066e-08, 
    6.473585e-08, 6.456669e-08, 6.519728e-08, 6.501806e-08, 6.553597e-08, 
    6.540572e-08, 6.552985e-08, 6.549221e-08, 6.553034e-08, 6.533932e-08, 
    6.542116e-08, 6.525307e-08, 6.459837e-08, 6.479079e-08, 6.421691e-08, 
    6.387185e-08, 6.364264e-08, 6.347999e-08, 6.350298e-08, 6.354682e-08, 
    6.377208e-08, 6.398385e-08, 6.414524e-08, 6.42532e-08, 6.435957e-08, 
    6.468156e-08, 6.485197e-08, 6.523354e-08, 6.516466e-08, 6.528133e-08, 
    6.539276e-08, 6.557987e-08, 6.554907e-08, 6.563151e-08, 6.527824e-08, 
    6.551303e-08, 6.512544e-08, 6.523145e-08, 6.438852e-08, 6.406734e-08, 
    6.393085e-08, 6.381136e-08, 6.352067e-08, 6.372141e-08, 6.364228e-08, 
    6.383054e-08, 6.395017e-08, 6.3891e-08, 6.425615e-08, 6.411419e-08, 
    6.486207e-08, 6.453993e-08, 6.537977e-08, 6.51788e-08, 6.542793e-08, 
    6.53008e-08, 6.551863e-08, 6.532259e-08, 6.566219e-08, 6.573613e-08, 
    6.56856e-08, 6.587971e-08, 6.531172e-08, 6.552985e-08, 6.388935e-08, 
    6.389899e-08, 6.394394e-08, 6.374634e-08, 6.373425e-08, 6.355315e-08, 
    6.371429e-08, 6.378291e-08, 6.39571e-08, 6.406013e-08, 6.415808e-08, 
    6.437342e-08, 6.461393e-08, 6.495023e-08, 6.519183e-08, 6.535377e-08, 
    6.525447e-08, 6.534214e-08, 6.524414e-08, 6.519819e-08, 6.570843e-08, 
    6.542193e-08, 6.585179e-08, 6.5828e-08, 6.563347e-08, 6.583068e-08, 
    6.390577e-08, 6.385024e-08, 6.365745e-08, 6.380832e-08, 6.353343e-08, 
    6.36873e-08, 6.377579e-08, 6.411717e-08, 6.419216e-08, 6.426171e-08, 
    6.439907e-08, 6.457535e-08, 6.488458e-08, 6.515364e-08, 6.539925e-08, 
    6.538125e-08, 6.538759e-08, 6.544246e-08, 6.530654e-08, 6.546477e-08, 
    6.549133e-08, 6.542189e-08, 6.582482e-08, 6.570971e-08, 6.58275e-08, 
    6.575254e-08, 6.386828e-08, 6.396172e-08, 6.391124e-08, 6.400618e-08, 
    6.393929e-08, 6.423671e-08, 6.432588e-08, 6.474312e-08, 6.457188e-08, 
    6.484441e-08, 6.459956e-08, 6.464295e-08, 6.485331e-08, 6.461279e-08, 
    6.513881e-08, 6.47822e-08, 6.544459e-08, 6.508849e-08, 6.546691e-08, 
    6.539818e-08, 6.551196e-08, 6.561386e-08, 6.574206e-08, 6.59786e-08, 
    6.592382e-08, 6.612164e-08, 6.410102e-08, 6.422221e-08, 6.421153e-08, 
    6.433836e-08, 6.443215e-08, 6.463544e-08, 6.496149e-08, 6.483888e-08, 
    6.506396e-08, 6.510916e-08, 6.476719e-08, 6.497716e-08, 6.430331e-08, 
    6.441219e-08, 6.434736e-08, 6.411058e-08, 6.486714e-08, 6.447888e-08, 
    6.519582e-08, 6.498549e-08, 6.559934e-08, 6.529407e-08, 6.589367e-08, 
    6.615002e-08, 6.639124e-08, 6.667317e-08, 6.428834e-08, 6.4206e-08, 
    6.435344e-08, 6.455743e-08, 6.47467e-08, 6.499832e-08, 6.502406e-08, 
    6.507121e-08, 6.51933e-08, 6.529596e-08, 6.508611e-08, 6.53217e-08, 
    6.443745e-08, 6.490084e-08, 6.417487e-08, 6.439348e-08, 6.454541e-08, 
    6.447876e-08, 6.482487e-08, 6.490644e-08, 6.523793e-08, 6.506657e-08, 
    6.608675e-08, 6.56354e-08, 6.688783e-08, 6.653783e-08, 6.417723e-08, 
    6.428806e-08, 6.467379e-08, 6.449026e-08, 6.501512e-08, 6.514431e-08, 
    6.524932e-08, 6.538358e-08, 6.539807e-08, 6.547761e-08, 6.534727e-08, 
    6.547247e-08, 6.499886e-08, 6.52105e-08, 6.46297e-08, 6.477106e-08, 
    6.470603e-08, 6.463469e-08, 6.485485e-08, 6.508942e-08, 6.509442e-08, 
    6.516963e-08, 6.53816e-08, 6.501724e-08, 6.614502e-08, 6.544855e-08, 
    6.440892e-08, 6.462241e-08, 6.465289e-08, 6.457019e-08, 6.513136e-08, 
    6.492802e-08, 6.547567e-08, 6.532767e-08, 6.557018e-08, 6.544967e-08, 
    6.543194e-08, 6.527716e-08, 6.51808e-08, 6.493735e-08, 6.473926e-08, 
    6.458218e-08, 6.46187e-08, 6.479126e-08, 6.510376e-08, 6.539939e-08, 
    6.533463e-08, 6.555175e-08, 6.497706e-08, 6.521804e-08, 6.512491e-08, 
    6.536776e-08, 6.483562e-08, 6.528879e-08, 6.471979e-08, 6.476968e-08, 
    6.492399e-08, 6.52344e-08, 6.530306e-08, 6.537638e-08, 6.533113e-08, 
    6.51117e-08, 6.507574e-08, 6.492024e-08, 6.487731e-08, 6.475882e-08, 
    6.466072e-08, 6.475035e-08, 6.484448e-08, 6.511178e-08, 6.535268e-08, 
    6.561532e-08, 6.567959e-08, 6.598647e-08, 6.573666e-08, 6.61489e-08, 
    6.579844e-08, 6.64051e-08, 6.531504e-08, 6.578811e-08, 6.493101e-08, 
    6.502334e-08, 6.519036e-08, 6.557342e-08, 6.536661e-08, 6.560847e-08, 
    6.507433e-08, 6.479721e-08, 6.47255e-08, 6.459173e-08, 6.472857e-08, 
    6.471743e-08, 6.484837e-08, 6.480629e-08, 6.512066e-08, 6.49518e-08, 
    6.54315e-08, 6.560656e-08, 6.610091e-08, 6.640397e-08, 6.671245e-08, 
    6.684864e-08, 6.689009e-08, 6.690742e-08 ;

 HR_vr =
  2.669659e-07, 2.676731e-07, 2.675357e-07, 2.681056e-07, 2.677895e-07, 
    2.681626e-07, 2.671093e-07, 2.677012e-07, 2.673234e-07, 2.670296e-07, 
    2.692103e-07, 2.68131e-07, 2.703289e-07, 2.696422e-07, 2.713656e-07, 
    2.702222e-07, 2.715959e-07, 2.713326e-07, 2.721245e-07, 2.718978e-07, 
    2.729097e-07, 2.722292e-07, 2.734334e-07, 2.727472e-07, 2.728546e-07, 
    2.722067e-07, 2.683483e-07, 2.69076e-07, 2.683052e-07, 2.68409e-07, 
    2.683624e-07, 2.677961e-07, 2.675105e-07, 2.669118e-07, 2.670205e-07, 
    2.674602e-07, 2.684557e-07, 2.681179e-07, 2.689687e-07, 2.689495e-07, 
    2.698954e-07, 2.694691e-07, 2.710565e-07, 2.706058e-07, 2.719072e-07, 
    2.715802e-07, 2.718919e-07, 2.717974e-07, 2.718931e-07, 2.714134e-07, 
    2.71619e-07, 2.711967e-07, 2.69549e-07, 2.700338e-07, 2.685868e-07, 
    2.677151e-07, 2.671353e-07, 2.667236e-07, 2.667818e-07, 2.668928e-07, 
    2.674628e-07, 2.679981e-07, 2.684058e-07, 2.686783e-07, 2.689468e-07, 
    2.697587e-07, 2.701878e-07, 2.711476e-07, 2.709744e-07, 2.712677e-07, 
    2.715476e-07, 2.720174e-07, 2.719401e-07, 2.72147e-07, 2.712599e-07, 
    2.718496e-07, 2.708759e-07, 2.711423e-07, 2.690199e-07, 2.68209e-07, 
    2.678642e-07, 2.675621e-07, 2.668266e-07, 2.673346e-07, 2.671344e-07, 
    2.676106e-07, 2.67913e-07, 2.677634e-07, 2.686858e-07, 2.683274e-07, 
    2.702132e-07, 2.694017e-07, 2.71515e-07, 2.7101e-07, 2.71636e-07, 
    2.713166e-07, 2.718637e-07, 2.713713e-07, 2.72224e-07, 2.724095e-07, 
    2.722827e-07, 2.727694e-07, 2.71344e-07, 2.718919e-07, 2.677592e-07, 
    2.677837e-07, 2.678973e-07, 2.673977e-07, 2.673671e-07, 2.669088e-07, 
    2.673166e-07, 2.674902e-07, 2.679305e-07, 2.681909e-07, 2.684382e-07, 
    2.689818e-07, 2.695882e-07, 2.704351e-07, 2.710427e-07, 2.714497e-07, 
    2.712002e-07, 2.714205e-07, 2.711742e-07, 2.710587e-07, 2.7234e-07, 
    2.716209e-07, 2.726995e-07, 2.726398e-07, 2.721519e-07, 2.726465e-07, 
    2.678008e-07, 2.676604e-07, 2.671728e-07, 2.675544e-07, 2.668589e-07, 
    2.672483e-07, 2.674722e-07, 2.683349e-07, 2.685243e-07, 2.686998e-07, 
    2.690464e-07, 2.694909e-07, 2.702699e-07, 2.709467e-07, 2.715639e-07, 
    2.715187e-07, 2.715346e-07, 2.716724e-07, 2.71331e-07, 2.717285e-07, 
    2.717952e-07, 2.716208e-07, 2.726318e-07, 2.723432e-07, 2.726385e-07, 
    2.724506e-07, 2.67706e-07, 2.679422e-07, 2.678146e-07, 2.680545e-07, 
    2.678855e-07, 2.686368e-07, 2.688618e-07, 2.699137e-07, 2.694822e-07, 
    2.701688e-07, 2.695519e-07, 2.696613e-07, 2.701912e-07, 2.695853e-07, 
    2.709095e-07, 2.700121e-07, 2.716778e-07, 2.70783e-07, 2.717338e-07, 
    2.715612e-07, 2.718469e-07, 2.721027e-07, 2.724243e-07, 2.730173e-07, 
    2.7288e-07, 2.733755e-07, 2.682941e-07, 2.686001e-07, 2.685732e-07, 
    2.688933e-07, 2.691299e-07, 2.696424e-07, 2.704634e-07, 2.701548e-07, 
    2.707212e-07, 2.708349e-07, 2.699743e-07, 2.705029e-07, 2.688049e-07, 
    2.690796e-07, 2.68916e-07, 2.683183e-07, 2.70226e-07, 2.692477e-07, 
    2.710528e-07, 2.705238e-07, 2.720663e-07, 2.712997e-07, 2.728044e-07, 
    2.734466e-07, 2.740501e-07, 2.747547e-07, 2.687671e-07, 2.685592e-07, 
    2.689313e-07, 2.694458e-07, 2.699227e-07, 2.705561e-07, 2.706209e-07, 
    2.707395e-07, 2.710464e-07, 2.713044e-07, 2.70777e-07, 2.713691e-07, 
    2.691433e-07, 2.703108e-07, 2.684806e-07, 2.690324e-07, 2.694155e-07, 
    2.692474e-07, 2.701195e-07, 2.703249e-07, 2.711586e-07, 2.707278e-07, 
    2.732882e-07, 2.721568e-07, 2.752905e-07, 2.744165e-07, 2.684866e-07, 
    2.687663e-07, 2.69739e-07, 2.692764e-07, 2.705983e-07, 2.709232e-07, 
    2.711872e-07, 2.715246e-07, 2.71561e-07, 2.717607e-07, 2.714334e-07, 
    2.717478e-07, 2.705575e-07, 2.710897e-07, 2.696279e-07, 2.69984e-07, 
    2.698202e-07, 2.696405e-07, 2.70195e-07, 2.707853e-07, 2.707978e-07, 
    2.709869e-07, 2.715198e-07, 2.706037e-07, 2.734342e-07, 2.716879e-07, 
    2.690713e-07, 2.696096e-07, 2.696863e-07, 2.694779e-07, 2.708908e-07, 
    2.703792e-07, 2.717559e-07, 2.713841e-07, 2.719931e-07, 2.716906e-07, 
    2.71646e-07, 2.712572e-07, 2.71015e-07, 2.704027e-07, 2.699039e-07, 
    2.695081e-07, 2.696002e-07, 2.700349e-07, 2.708214e-07, 2.715643e-07, 
    2.714016e-07, 2.719468e-07, 2.705026e-07, 2.711086e-07, 2.708745e-07, 
    2.714848e-07, 2.701466e-07, 2.712866e-07, 2.698549e-07, 2.699805e-07, 
    2.703691e-07, 2.711498e-07, 2.713223e-07, 2.715065e-07, 2.713928e-07, 
    2.708413e-07, 2.707509e-07, 2.703596e-07, 2.702516e-07, 2.699532e-07, 
    2.69706e-07, 2.699319e-07, 2.701689e-07, 2.708415e-07, 2.71447e-07, 
    2.721064e-07, 2.722676e-07, 2.73037e-07, 2.724109e-07, 2.734439e-07, 
    2.725658e-07, 2.740848e-07, 2.713524e-07, 2.725399e-07, 2.703867e-07, 
    2.706191e-07, 2.710391e-07, 2.720013e-07, 2.71482e-07, 2.720892e-07, 
    2.707473e-07, 2.700499e-07, 2.698693e-07, 2.695322e-07, 2.69877e-07, 
    2.69849e-07, 2.701787e-07, 2.700727e-07, 2.708638e-07, 2.70439e-07, 
    2.716449e-07, 2.720844e-07, 2.733236e-07, 2.740819e-07, 2.748527e-07, 
    2.751927e-07, 2.752961e-07, 2.753393e-07,
  2.414858e-07, 2.423968e-07, 2.422197e-07, 2.42954e-07, 2.425468e-07, 
    2.430274e-07, 2.416706e-07, 2.424329e-07, 2.419463e-07, 2.415678e-07, 
    2.443772e-07, 2.429867e-07, 2.458195e-07, 2.449343e-07, 2.471562e-07, 
    2.456817e-07, 2.474533e-07, 2.471138e-07, 2.481353e-07, 2.478427e-07, 
    2.491479e-07, 2.482702e-07, 2.498238e-07, 2.489384e-07, 2.49077e-07, 
    2.482413e-07, 2.432668e-07, 2.442042e-07, 2.432112e-07, 2.433449e-07, 
    2.432849e-07, 2.425552e-07, 2.421872e-07, 2.414161e-07, 2.415562e-07, 
    2.421225e-07, 2.434051e-07, 2.429699e-07, 2.440663e-07, 2.440416e-07, 
    2.452606e-07, 2.447112e-07, 2.467577e-07, 2.461765e-07, 2.47855e-07, 
    2.474331e-07, 2.478351e-07, 2.477133e-07, 2.478367e-07, 2.47218e-07, 
    2.474831e-07, 2.469385e-07, 2.448141e-07, 2.45439e-07, 2.43574e-07, 
    2.424507e-07, 2.41704e-07, 2.411737e-07, 2.412487e-07, 2.413916e-07, 
    2.421258e-07, 2.428156e-07, 2.433408e-07, 2.436921e-07, 2.44038e-07, 
    2.450842e-07, 2.456375e-07, 2.468751e-07, 2.46652e-07, 2.4703e-07, 
    2.473912e-07, 2.479971e-07, 2.478974e-07, 2.481642e-07, 2.470201e-07, 
    2.477806e-07, 2.465248e-07, 2.468684e-07, 2.441319e-07, 2.430873e-07, 
    2.426429e-07, 2.422538e-07, 2.413063e-07, 2.419607e-07, 2.417028e-07, 
    2.423163e-07, 2.427059e-07, 2.425132e-07, 2.437017e-07, 2.432398e-07, 
    2.456703e-07, 2.446242e-07, 2.47349e-07, 2.466978e-07, 2.475051e-07, 
    2.470932e-07, 2.477988e-07, 2.471638e-07, 2.482635e-07, 2.485028e-07, 
    2.483393e-07, 2.489672e-07, 2.471286e-07, 2.478351e-07, 2.425078e-07, 
    2.425392e-07, 2.426856e-07, 2.420419e-07, 2.420026e-07, 2.414123e-07, 
    2.419375e-07, 2.421611e-07, 2.427285e-07, 2.430639e-07, 2.433826e-07, 
    2.44083e-07, 2.448646e-07, 2.459564e-07, 2.4674e-07, 2.472649e-07, 
    2.469431e-07, 2.472272e-07, 2.469096e-07, 2.467607e-07, 2.484131e-07, 
    2.474856e-07, 2.488769e-07, 2.488e-07, 2.481706e-07, 2.488086e-07, 
    2.425613e-07, 2.423805e-07, 2.417523e-07, 2.422439e-07, 2.41348e-07, 
    2.418496e-07, 2.421378e-07, 2.432494e-07, 2.434935e-07, 2.437197e-07, 
    2.441664e-07, 2.447393e-07, 2.457434e-07, 2.466162e-07, 2.474122e-07, 
    2.473539e-07, 2.473744e-07, 2.475521e-07, 2.471118e-07, 2.476244e-07, 
    2.477104e-07, 2.474855e-07, 2.487897e-07, 2.484173e-07, 2.487984e-07, 
    2.485559e-07, 2.424393e-07, 2.427435e-07, 2.425791e-07, 2.428882e-07, 
    2.426704e-07, 2.436384e-07, 2.439284e-07, 2.452842e-07, 2.44728e-07, 
    2.45613e-07, 2.44818e-07, 2.449589e-07, 2.456418e-07, 2.44861e-07, 
    2.46568e-07, 2.45411e-07, 2.47559e-07, 2.464049e-07, 2.476313e-07, 
    2.474087e-07, 2.477772e-07, 2.481071e-07, 2.48522e-07, 2.492869e-07, 
    2.491098e-07, 2.497491e-07, 2.431969e-07, 2.435912e-07, 2.435565e-07, 
    2.43969e-07, 2.442739e-07, 2.449345e-07, 2.45993e-07, 2.455951e-07, 
    2.463254e-07, 2.46472e-07, 2.453624e-07, 2.460438e-07, 2.43855e-07, 
    2.44209e-07, 2.439983e-07, 2.43228e-07, 2.456868e-07, 2.444258e-07, 
    2.467529e-07, 2.460709e-07, 2.480601e-07, 2.470713e-07, 2.490123e-07, 
    2.498407e-07, 2.506197e-07, 2.51529e-07, 2.438064e-07, 2.435385e-07, 
    2.440181e-07, 2.44681e-07, 2.452958e-07, 2.461125e-07, 2.46196e-07, 
    2.463489e-07, 2.467448e-07, 2.470775e-07, 2.463972e-07, 2.471609e-07, 
    2.44291e-07, 2.457962e-07, 2.434372e-07, 2.441482e-07, 2.44642e-07, 
    2.444254e-07, 2.455496e-07, 2.458144e-07, 2.468894e-07, 2.463339e-07, 
    2.496363e-07, 2.481767e-07, 2.522208e-07, 2.510926e-07, 2.434449e-07, 
    2.438055e-07, 2.450591e-07, 2.444628e-07, 2.46167e-07, 2.465859e-07, 
    2.469264e-07, 2.473614e-07, 2.474084e-07, 2.47666e-07, 2.472438e-07, 
    2.476493e-07, 2.461142e-07, 2.468005e-07, 2.449159e-07, 2.45375e-07, 
    2.451638e-07, 2.449321e-07, 2.45647e-07, 2.464079e-07, 2.464242e-07, 
    2.46668e-07, 2.473548e-07, 2.461739e-07, 2.498244e-07, 2.475716e-07, 
    2.441984e-07, 2.448921e-07, 2.449912e-07, 2.447225e-07, 2.46544e-07, 
    2.458844e-07, 2.476597e-07, 2.471803e-07, 2.479657e-07, 2.475755e-07, 
    2.475181e-07, 2.470166e-07, 2.467042e-07, 2.459147e-07, 2.452717e-07, 
    2.447615e-07, 2.448802e-07, 2.454405e-07, 2.464544e-07, 2.474126e-07, 
    2.472028e-07, 2.479061e-07, 2.460435e-07, 2.46825e-07, 2.46523e-07, 
    2.473101e-07, 2.455845e-07, 2.470541e-07, 2.452085e-07, 2.453705e-07, 
    2.458713e-07, 2.468779e-07, 2.471005e-07, 2.473381e-07, 2.471915e-07, 
    2.464802e-07, 2.463636e-07, 2.458592e-07, 2.457198e-07, 2.453352e-07, 
    2.450167e-07, 2.453077e-07, 2.456133e-07, 2.464805e-07, 2.472613e-07, 
    2.481118e-07, 2.483198e-07, 2.493122e-07, 2.485044e-07, 2.49837e-07, 
    2.487041e-07, 2.506642e-07, 2.471392e-07, 2.486708e-07, 2.458941e-07, 
    2.461937e-07, 2.467352e-07, 2.479761e-07, 2.473064e-07, 2.480896e-07, 
    2.46359e-07, 2.454598e-07, 2.452271e-07, 2.447925e-07, 2.45237e-07, 
    2.452008e-07, 2.456259e-07, 2.454894e-07, 2.465093e-07, 2.459616e-07, 
    2.475166e-07, 2.480834e-07, 2.496821e-07, 2.506607e-07, 2.516557e-07, 
    2.520946e-07, 2.522281e-07, 2.522839e-07,
  2.259477e-07, 2.26945e-07, 2.267512e-07, 2.275552e-07, 2.271093e-07, 
    2.276357e-07, 2.2615e-07, 2.269846e-07, 2.264519e-07, 2.260376e-07, 
    2.291142e-07, 2.275911e-07, 2.306949e-07, 2.297247e-07, 2.321607e-07, 
    2.305439e-07, 2.324865e-07, 2.321141e-07, 2.332346e-07, 2.329137e-07, 
    2.343459e-07, 2.333827e-07, 2.350877e-07, 2.341159e-07, 2.34268e-07, 
    2.333509e-07, 2.278978e-07, 2.289247e-07, 2.278369e-07, 2.279834e-07, 
    2.279177e-07, 2.271185e-07, 2.267156e-07, 2.258715e-07, 2.260248e-07, 
    2.266447e-07, 2.280493e-07, 2.275727e-07, 2.287736e-07, 2.287465e-07, 
    2.300823e-07, 2.294802e-07, 2.317236e-07, 2.310863e-07, 2.329271e-07, 
    2.324644e-07, 2.329054e-07, 2.327717e-07, 2.329071e-07, 2.322284e-07, 
    2.325192e-07, 2.319219e-07, 2.29593e-07, 2.302778e-07, 2.282343e-07, 
    2.270041e-07, 2.261866e-07, 2.256062e-07, 2.256882e-07, 2.258447e-07, 
    2.266484e-07, 2.274036e-07, 2.279789e-07, 2.283636e-07, 2.287426e-07, 
    2.29889e-07, 2.304955e-07, 2.318524e-07, 2.316076e-07, 2.320223e-07, 
    2.324183e-07, 2.33083e-07, 2.329736e-07, 2.332664e-07, 2.320114e-07, 
    2.328456e-07, 2.314682e-07, 2.31845e-07, 2.288455e-07, 2.277012e-07, 
    2.272145e-07, 2.267885e-07, 2.257513e-07, 2.264676e-07, 2.261853e-07, 
    2.268569e-07, 2.272835e-07, 2.270725e-07, 2.283741e-07, 2.278683e-07, 
    2.305314e-07, 2.293849e-07, 2.323722e-07, 2.316579e-07, 2.325433e-07, 
    2.320916e-07, 2.328655e-07, 2.32169e-07, 2.333753e-07, 2.336378e-07, 
    2.334585e-07, 2.341475e-07, 2.321304e-07, 2.329054e-07, 2.270666e-07, 
    2.27101e-07, 2.272614e-07, 2.265566e-07, 2.265134e-07, 2.258673e-07, 
    2.264423e-07, 2.26687e-07, 2.273082e-07, 2.276756e-07, 2.280247e-07, 
    2.287919e-07, 2.296483e-07, 2.30845e-07, 2.317042e-07, 2.322798e-07, 
    2.319269e-07, 2.322385e-07, 2.318902e-07, 2.317269e-07, 2.335395e-07, 
    2.325219e-07, 2.340484e-07, 2.33964e-07, 2.332733e-07, 2.339735e-07, 
    2.271252e-07, 2.269272e-07, 2.262394e-07, 2.267777e-07, 2.257969e-07, 
    2.26346e-07, 2.266616e-07, 2.278788e-07, 2.281461e-07, 2.283939e-07, 
    2.288833e-07, 2.29511e-07, 2.306115e-07, 2.315684e-07, 2.324414e-07, 
    2.323774e-07, 2.324e-07, 2.325949e-07, 2.32112e-07, 2.326742e-07, 
    2.327685e-07, 2.325218e-07, 2.339527e-07, 2.335441e-07, 2.339622e-07, 
    2.336962e-07, 2.269916e-07, 2.273247e-07, 2.271447e-07, 2.274832e-07, 
    2.272447e-07, 2.283048e-07, 2.286225e-07, 2.301081e-07, 2.294986e-07, 
    2.304686e-07, 2.295972e-07, 2.297516e-07, 2.305001e-07, 2.296443e-07, 
    2.315156e-07, 2.302472e-07, 2.326025e-07, 2.313367e-07, 2.326818e-07, 
    2.324376e-07, 2.328418e-07, 2.332037e-07, 2.336589e-07, 2.344984e-07, 
    2.34304e-07, 2.350058e-07, 2.278213e-07, 2.282532e-07, 2.282152e-07, 
    2.28667e-07, 2.290011e-07, 2.297249e-07, 2.308851e-07, 2.30449e-07, 
    2.312496e-07, 2.314103e-07, 2.301939e-07, 2.309408e-07, 2.285421e-07, 
    2.289299e-07, 2.286991e-07, 2.278554e-07, 2.305494e-07, 2.291674e-07, 
    2.317184e-07, 2.309705e-07, 2.331521e-07, 2.320675e-07, 2.34197e-07, 
    2.351063e-07, 2.359616e-07, 2.369604e-07, 2.284888e-07, 2.281954e-07, 
    2.287208e-07, 2.294472e-07, 2.301209e-07, 2.310161e-07, 2.311077e-07, 
    2.312753e-07, 2.317094e-07, 2.320744e-07, 2.313283e-07, 2.321658e-07, 
    2.290198e-07, 2.306694e-07, 2.280845e-07, 2.288633e-07, 2.294044e-07, 
    2.291671e-07, 2.303991e-07, 2.306893e-07, 2.31868e-07, 2.312589e-07, 
    2.348819e-07, 2.332801e-07, 2.377204e-07, 2.36481e-07, 2.280929e-07, 
    2.284878e-07, 2.298614e-07, 2.29208e-07, 2.310759e-07, 2.315353e-07, 
    2.319086e-07, 2.323857e-07, 2.324372e-07, 2.327198e-07, 2.322567e-07, 
    2.327015e-07, 2.31018e-07, 2.317706e-07, 2.297045e-07, 2.302076e-07, 
    2.299762e-07, 2.297223e-07, 2.305058e-07, 2.313401e-07, 2.313579e-07, 
    2.316253e-07, 2.323784e-07, 2.310834e-07, 2.350885e-07, 2.326163e-07, 
    2.289184e-07, 2.296784e-07, 2.29787e-07, 2.294926e-07, 2.314892e-07, 
    2.307661e-07, 2.327129e-07, 2.32187e-07, 2.330486e-07, 2.326205e-07, 
    2.325575e-07, 2.320076e-07, 2.31665e-07, 2.307993e-07, 2.300945e-07, 
    2.295353e-07, 2.296654e-07, 2.302795e-07, 2.313911e-07, 2.324419e-07, 
    2.322117e-07, 2.329831e-07, 2.309405e-07, 2.317974e-07, 2.314662e-07, 
    2.323295e-07, 2.304374e-07, 2.320487e-07, 2.300252e-07, 2.302027e-07, 
    2.307517e-07, 2.318554e-07, 2.320996e-07, 2.323601e-07, 2.321994e-07, 
    2.314193e-07, 2.312915e-07, 2.307384e-07, 2.305857e-07, 2.301641e-07, 
    2.298149e-07, 2.301339e-07, 2.304688e-07, 2.314196e-07, 2.322759e-07, 
    2.332089e-07, 2.334371e-07, 2.345262e-07, 2.336396e-07, 2.351022e-07, 
    2.338588e-07, 2.360105e-07, 2.32142e-07, 2.338223e-07, 2.307767e-07, 
    2.311052e-07, 2.316989e-07, 2.3306e-07, 2.323254e-07, 2.331845e-07, 
    2.312864e-07, 2.303007e-07, 2.300455e-07, 2.295693e-07, 2.300564e-07, 
    2.300168e-07, 2.304827e-07, 2.30333e-07, 2.314512e-07, 2.308507e-07, 
    2.325559e-07, 2.331777e-07, 2.349322e-07, 2.360066e-07, 2.370995e-07, 
    2.375817e-07, 2.377284e-07, 2.377897e-07,
  2.166374e-07, 2.176639e-07, 2.174644e-07, 2.182922e-07, 2.17833e-07, 
    2.18375e-07, 2.168455e-07, 2.177047e-07, 2.171562e-07, 2.167298e-07, 
    2.198984e-07, 2.183291e-07, 2.21528e-07, 2.205275e-07, 2.230404e-07, 
    2.213723e-07, 2.233767e-07, 2.229923e-07, 2.241491e-07, 2.238177e-07, 
    2.252972e-07, 2.243021e-07, 2.260639e-07, 2.250596e-07, 2.252167e-07, 
    2.242692e-07, 2.18645e-07, 2.197031e-07, 2.185823e-07, 2.187332e-07, 
    2.186655e-07, 2.178425e-07, 2.174277e-07, 2.165589e-07, 2.167167e-07, 
    2.173548e-07, 2.18801e-07, 2.183101e-07, 2.195472e-07, 2.195193e-07, 
    2.208962e-07, 2.202755e-07, 2.225893e-07, 2.219317e-07, 2.238316e-07, 
    2.233539e-07, 2.238091e-07, 2.236711e-07, 2.238109e-07, 2.231103e-07, 
    2.234105e-07, 2.227939e-07, 2.203917e-07, 2.210978e-07, 2.189916e-07, 
    2.177248e-07, 2.168832e-07, 2.162859e-07, 2.163704e-07, 2.165313e-07, 
    2.173585e-07, 2.181361e-07, 2.187285e-07, 2.191248e-07, 2.195153e-07, 
    2.20697e-07, 2.213223e-07, 2.227222e-07, 2.224696e-07, 2.228975e-07, 
    2.233063e-07, 2.239926e-07, 2.238796e-07, 2.241819e-07, 2.228862e-07, 
    2.237474e-07, 2.223257e-07, 2.227146e-07, 2.196215e-07, 2.184426e-07, 
    2.179414e-07, 2.175027e-07, 2.164353e-07, 2.171725e-07, 2.168819e-07, 
    2.175732e-07, 2.180124e-07, 2.177951e-07, 2.191357e-07, 2.186145e-07, 
    2.213594e-07, 2.201773e-07, 2.232586e-07, 2.225215e-07, 2.234353e-07, 
    2.22969e-07, 2.23768e-07, 2.230489e-07, 2.242945e-07, 2.245656e-07, 
    2.243803e-07, 2.250921e-07, 2.230091e-07, 2.238091e-07, 2.177891e-07, 
    2.178245e-07, 2.179895e-07, 2.17264e-07, 2.172196e-07, 2.165546e-07, 
    2.171463e-07, 2.173983e-07, 2.180378e-07, 2.184161e-07, 2.187757e-07, 
    2.195661e-07, 2.204488e-07, 2.216829e-07, 2.225692e-07, 2.231633e-07, 
    2.22799e-07, 2.231207e-07, 2.227611e-07, 2.225926e-07, 2.24464e-07, 
    2.234133e-07, 2.249898e-07, 2.249025e-07, 2.241891e-07, 2.249124e-07, 
    2.178494e-07, 2.176455e-07, 2.169376e-07, 2.174916e-07, 2.164822e-07, 
    2.170472e-07, 2.173721e-07, 2.186254e-07, 2.189008e-07, 2.191561e-07, 
    2.196603e-07, 2.203072e-07, 2.21442e-07, 2.224291e-07, 2.233301e-07, 
    2.232641e-07, 2.232873e-07, 2.234886e-07, 2.229901e-07, 2.235704e-07, 
    2.236678e-07, 2.234132e-07, 2.248909e-07, 2.244687e-07, 2.249007e-07, 
    2.246258e-07, 2.177118e-07, 2.180548e-07, 2.178694e-07, 2.18218e-07, 
    2.179725e-07, 2.190643e-07, 2.193916e-07, 2.209229e-07, 2.202945e-07, 
    2.212946e-07, 2.203961e-07, 2.205553e-07, 2.213272e-07, 2.204446e-07, 
    2.223747e-07, 2.210663e-07, 2.234964e-07, 2.221901e-07, 2.235783e-07, 
    2.233262e-07, 2.237435e-07, 2.241172e-07, 2.245874e-07, 2.254547e-07, 
    2.252539e-07, 2.259792e-07, 2.185662e-07, 2.190111e-07, 2.189719e-07, 
    2.194374e-07, 2.197817e-07, 2.205278e-07, 2.217242e-07, 2.212743e-07, 
    2.221002e-07, 2.222659e-07, 2.210112e-07, 2.217816e-07, 2.193088e-07, 
    2.197084e-07, 2.194705e-07, 2.186013e-07, 2.21378e-07, 2.199532e-07, 
    2.225839e-07, 2.218122e-07, 2.24064e-07, 2.229443e-07, 2.251433e-07, 
    2.260831e-07, 2.269675e-07, 2.280007e-07, 2.192538e-07, 2.189516e-07, 
    2.194928e-07, 2.202415e-07, 2.20936e-07, 2.218593e-07, 2.219538e-07, 
    2.221267e-07, 2.225746e-07, 2.229512e-07, 2.221814e-07, 2.230456e-07, 
    2.198011e-07, 2.215016e-07, 2.188373e-07, 2.196397e-07, 2.201973e-07, 
    2.199527e-07, 2.212229e-07, 2.215222e-07, 2.227383e-07, 2.221097e-07, 
    2.258512e-07, 2.241962e-07, 2.287873e-07, 2.275047e-07, 2.18846e-07, 
    2.192528e-07, 2.206685e-07, 2.199949e-07, 2.219209e-07, 2.223949e-07, 
    2.227802e-07, 2.232726e-07, 2.233258e-07, 2.236175e-07, 2.231395e-07, 
    2.235987e-07, 2.218613e-07, 2.226377e-07, 2.205067e-07, 2.210254e-07, 
    2.207868e-07, 2.20525e-07, 2.213329e-07, 2.221935e-07, 2.222119e-07, 
    2.224878e-07, 2.232653e-07, 2.219287e-07, 2.260648e-07, 2.235109e-07, 
    2.196964e-07, 2.204799e-07, 2.205918e-07, 2.202883e-07, 2.223474e-07, 
    2.216014e-07, 2.236104e-07, 2.230675e-07, 2.23957e-07, 2.23515e-07, 
    2.2345e-07, 2.228823e-07, 2.225288e-07, 2.216356e-07, 2.209087e-07, 
    2.203323e-07, 2.204663e-07, 2.210995e-07, 2.222461e-07, 2.233306e-07, 
    2.230931e-07, 2.238894e-07, 2.217813e-07, 2.226654e-07, 2.223237e-07, 
    2.232146e-07, 2.212623e-07, 2.229249e-07, 2.208373e-07, 2.210204e-07, 
    2.215866e-07, 2.227254e-07, 2.229772e-07, 2.232462e-07, 2.230802e-07, 
    2.222752e-07, 2.221433e-07, 2.215728e-07, 2.214153e-07, 2.209805e-07, 
    2.206205e-07, 2.209494e-07, 2.212948e-07, 2.222756e-07, 2.231593e-07, 
    2.241226e-07, 2.243583e-07, 2.254835e-07, 2.245676e-07, 2.26079e-07, 
    2.247941e-07, 2.270182e-07, 2.230212e-07, 2.247562e-07, 2.216123e-07, 
    2.219511e-07, 2.225639e-07, 2.239689e-07, 2.232104e-07, 2.240974e-07, 
    2.221382e-07, 2.211214e-07, 2.208583e-07, 2.203674e-07, 2.208695e-07, 
    2.208287e-07, 2.213091e-07, 2.211547e-07, 2.223081e-07, 2.216886e-07, 
    2.234484e-07, 2.240904e-07, 2.259032e-07, 2.270141e-07, 2.281447e-07, 
    2.286437e-07, 2.287956e-07, 2.288591e-07,
  2.081373e-07, 2.091061e-07, 2.089177e-07, 2.096995e-07, 2.092658e-07, 
    2.097778e-07, 2.083337e-07, 2.091446e-07, 2.086269e-07, 2.082245e-07, 
    2.11218e-07, 2.097344e-07, 2.127605e-07, 2.118131e-07, 2.141941e-07, 
    2.126131e-07, 2.145131e-07, 2.141484e-07, 2.152462e-07, 2.149316e-07, 
    2.163369e-07, 2.153914e-07, 2.170658e-07, 2.16111e-07, 2.162603e-07, 
    2.153602e-07, 2.100328e-07, 2.110333e-07, 2.099735e-07, 2.101162e-07, 
    2.100521e-07, 2.092748e-07, 2.088832e-07, 2.080633e-07, 2.082121e-07, 
    2.088143e-07, 2.101803e-07, 2.097164e-07, 2.108857e-07, 2.108593e-07, 
    2.121622e-07, 2.115746e-07, 2.137662e-07, 2.131429e-07, 2.149447e-07, 
    2.144914e-07, 2.149234e-07, 2.147924e-07, 2.149252e-07, 2.142603e-07, 
    2.145451e-07, 2.139602e-07, 2.116846e-07, 2.12353e-07, 2.103604e-07, 
    2.091637e-07, 2.083692e-07, 2.078058e-07, 2.078854e-07, 2.080373e-07, 
    2.088178e-07, 2.09552e-07, 2.101117e-07, 2.104863e-07, 2.108555e-07, 
    2.119736e-07, 2.125657e-07, 2.138923e-07, 2.136527e-07, 2.140586e-07, 
    2.144463e-07, 2.150976e-07, 2.149904e-07, 2.152774e-07, 2.140478e-07, 
    2.148649e-07, 2.135163e-07, 2.13885e-07, 2.109561e-07, 2.098415e-07, 
    2.093683e-07, 2.089539e-07, 2.079467e-07, 2.086422e-07, 2.08368e-07, 
    2.090204e-07, 2.094352e-07, 2.0923e-07, 2.104966e-07, 2.10004e-07, 
    2.126008e-07, 2.114817e-07, 2.144011e-07, 2.137019e-07, 2.145687e-07, 
    2.141263e-07, 2.148844e-07, 2.142021e-07, 2.153842e-07, 2.156418e-07, 
    2.154658e-07, 2.161419e-07, 2.141643e-07, 2.149235e-07, 2.092243e-07, 
    2.092577e-07, 2.094136e-07, 2.087286e-07, 2.086867e-07, 2.080592e-07, 
    2.086175e-07, 2.088554e-07, 2.094592e-07, 2.098165e-07, 2.101563e-07, 
    2.109036e-07, 2.117387e-07, 2.129072e-07, 2.137472e-07, 2.143106e-07, 
    2.139651e-07, 2.142701e-07, 2.139292e-07, 2.137694e-07, 2.155453e-07, 
    2.145478e-07, 2.160447e-07, 2.159618e-07, 2.152842e-07, 2.159711e-07, 
    2.092812e-07, 2.090887e-07, 2.084205e-07, 2.089434e-07, 2.079909e-07, 
    2.08524e-07, 2.088307e-07, 2.100144e-07, 2.102745e-07, 2.105159e-07, 
    2.109926e-07, 2.116046e-07, 2.12679e-07, 2.136144e-07, 2.144688e-07, 
    2.144062e-07, 2.144283e-07, 2.146192e-07, 2.141463e-07, 2.146969e-07, 
    2.147894e-07, 2.145477e-07, 2.159507e-07, 2.155497e-07, 2.1596e-07, 
    2.156989e-07, 2.091513e-07, 2.094752e-07, 2.093002e-07, 2.096294e-07, 
    2.093975e-07, 2.104291e-07, 2.107386e-07, 2.121874e-07, 2.115926e-07, 
    2.125394e-07, 2.116887e-07, 2.118394e-07, 2.125704e-07, 2.117347e-07, 
    2.135629e-07, 2.123232e-07, 2.146267e-07, 2.133879e-07, 2.147043e-07, 
    2.144651e-07, 2.148611e-07, 2.152159e-07, 2.156624e-07, 2.164866e-07, 
    2.162957e-07, 2.169852e-07, 2.099583e-07, 2.103788e-07, 2.103417e-07, 
    2.107818e-07, 2.111074e-07, 2.118133e-07, 2.129463e-07, 2.125201e-07, 
    2.133025e-07, 2.134597e-07, 2.12271e-07, 2.130008e-07, 2.106602e-07, 
    2.110382e-07, 2.108131e-07, 2.099915e-07, 2.126184e-07, 2.112697e-07, 
    2.137611e-07, 2.130297e-07, 2.151654e-07, 2.141029e-07, 2.161906e-07, 
    2.170842e-07, 2.179255e-07, 2.189097e-07, 2.106083e-07, 2.103225e-07, 
    2.108342e-07, 2.115425e-07, 2.121998e-07, 2.130743e-07, 2.131638e-07, 
    2.133277e-07, 2.137523e-07, 2.141094e-07, 2.133796e-07, 2.14199e-07, 
    2.111259e-07, 2.127355e-07, 2.102146e-07, 2.109732e-07, 2.115007e-07, 
    2.112692e-07, 2.124714e-07, 2.127549e-07, 2.139076e-07, 2.133116e-07, 
    2.168636e-07, 2.15291e-07, 2.196594e-07, 2.184372e-07, 2.102227e-07, 
    2.106073e-07, 2.119466e-07, 2.113092e-07, 2.131327e-07, 2.135819e-07, 
    2.139472e-07, 2.144144e-07, 2.144648e-07, 2.147416e-07, 2.14288e-07, 
    2.147237e-07, 2.130762e-07, 2.138122e-07, 2.117934e-07, 2.122845e-07, 
    2.120585e-07, 2.118107e-07, 2.125756e-07, 2.133911e-07, 2.134084e-07, 
    2.1367e-07, 2.144076e-07, 2.131401e-07, 2.170669e-07, 2.146406e-07, 
    2.110267e-07, 2.117681e-07, 2.118739e-07, 2.115867e-07, 2.135369e-07, 
    2.1283e-07, 2.147349e-07, 2.142198e-07, 2.150638e-07, 2.146443e-07, 
    2.145826e-07, 2.140441e-07, 2.137089e-07, 2.128624e-07, 2.12174e-07, 
    2.116283e-07, 2.117552e-07, 2.123547e-07, 2.13441e-07, 2.144694e-07, 
    2.14244e-07, 2.149997e-07, 2.130004e-07, 2.138384e-07, 2.135145e-07, 
    2.143593e-07, 2.125088e-07, 2.140847e-07, 2.121063e-07, 2.122797e-07, 
    2.128159e-07, 2.138953e-07, 2.141341e-07, 2.143893e-07, 2.142318e-07, 
    2.134685e-07, 2.133435e-07, 2.128029e-07, 2.126537e-07, 2.122419e-07, 
    2.119011e-07, 2.122125e-07, 2.125396e-07, 2.134688e-07, 2.143068e-07, 
    2.15221e-07, 2.154448e-07, 2.165141e-07, 2.156437e-07, 2.170804e-07, 
    2.15859e-07, 2.17974e-07, 2.141759e-07, 2.158229e-07, 2.128403e-07, 
    2.131613e-07, 2.137422e-07, 2.150752e-07, 2.143553e-07, 2.151972e-07, 
    2.133386e-07, 2.123754e-07, 2.121262e-07, 2.116615e-07, 2.121368e-07, 
    2.120981e-07, 2.125531e-07, 2.124069e-07, 2.134997e-07, 2.129126e-07, 
    2.145811e-07, 2.151905e-07, 2.169129e-07, 2.1797e-07, 2.190467e-07, 
    2.195224e-07, 2.196672e-07, 2.197278e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HTOP =
  0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823 ;

 INT_SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAISHA =
  0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503 ;

 LAISUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAKEICEFRAC =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAKEICETHICK =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAND_UPTAKE =
  6.35757e-08, 6.385525e-08, 6.38009e-08, 6.402639e-08, 6.39013e-08, 
    6.404895e-08, 6.363237e-08, 6.386636e-08, 6.371699e-08, 6.360087e-08, 
    6.446398e-08, 6.403645e-08, 6.490803e-08, 6.463537e-08, 6.532027e-08, 
    6.48656e-08, 6.541195e-08, 6.530715e-08, 6.562256e-08, 6.55322e-08, 
    6.593564e-08, 6.566426e-08, 6.614476e-08, 6.587083e-08, 6.591368e-08, 
    6.565531e-08, 6.412248e-08, 6.441076e-08, 6.41054e-08, 6.41465e-08, 
    6.412806e-08, 6.390389e-08, 6.379094e-08, 6.355432e-08, 6.359728e-08, 
    6.377105e-08, 6.416499e-08, 6.403126e-08, 6.436827e-08, 6.436066e-08, 
    6.473585e-08, 6.456669e-08, 6.519728e-08, 6.501806e-08, 6.553597e-08, 
    6.540572e-08, 6.552985e-08, 6.549221e-08, 6.553034e-08, 6.533932e-08, 
    6.542116e-08, 6.525307e-08, 6.459837e-08, 6.479079e-08, 6.421691e-08, 
    6.387185e-08, 6.364264e-08, 6.347999e-08, 6.350298e-08, 6.354682e-08, 
    6.377208e-08, 6.398385e-08, 6.414524e-08, 6.42532e-08, 6.435957e-08, 
    6.468156e-08, 6.485197e-08, 6.523354e-08, 6.516466e-08, 6.528133e-08, 
    6.539276e-08, 6.557987e-08, 6.554907e-08, 6.563151e-08, 6.527824e-08, 
    6.551303e-08, 6.512544e-08, 6.523145e-08, 6.438852e-08, 6.406734e-08, 
    6.393085e-08, 6.381136e-08, 6.352067e-08, 6.372141e-08, 6.364228e-08, 
    6.383054e-08, 6.395017e-08, 6.3891e-08, 6.425615e-08, 6.411419e-08, 
    6.486207e-08, 6.453993e-08, 6.537977e-08, 6.51788e-08, 6.542793e-08, 
    6.53008e-08, 6.551863e-08, 6.532259e-08, 6.566219e-08, 6.573613e-08, 
    6.56856e-08, 6.587971e-08, 6.531172e-08, 6.552985e-08, 6.388935e-08, 
    6.389899e-08, 6.394394e-08, 6.374634e-08, 6.373425e-08, 6.355315e-08, 
    6.371429e-08, 6.378291e-08, 6.39571e-08, 6.406013e-08, 6.415808e-08, 
    6.437342e-08, 6.461393e-08, 6.495023e-08, 6.519183e-08, 6.535377e-08, 
    6.525447e-08, 6.534214e-08, 6.524414e-08, 6.519819e-08, 6.570843e-08, 
    6.542193e-08, 6.585179e-08, 6.5828e-08, 6.563347e-08, 6.583068e-08, 
    6.390577e-08, 6.385024e-08, 6.365745e-08, 6.380832e-08, 6.353343e-08, 
    6.36873e-08, 6.377579e-08, 6.411717e-08, 6.419216e-08, 6.426171e-08, 
    6.439907e-08, 6.457535e-08, 6.488458e-08, 6.515364e-08, 6.539925e-08, 
    6.538125e-08, 6.538759e-08, 6.544246e-08, 6.530654e-08, 6.546477e-08, 
    6.549133e-08, 6.542189e-08, 6.582482e-08, 6.570971e-08, 6.58275e-08, 
    6.575254e-08, 6.386828e-08, 6.396172e-08, 6.391124e-08, 6.400618e-08, 
    6.393929e-08, 6.423671e-08, 6.432588e-08, 6.474312e-08, 6.457188e-08, 
    6.484441e-08, 6.459956e-08, 6.464295e-08, 6.485331e-08, 6.461279e-08, 
    6.513881e-08, 6.47822e-08, 6.544459e-08, 6.508849e-08, 6.546691e-08, 
    6.539818e-08, 6.551196e-08, 6.561386e-08, 6.574206e-08, 6.59786e-08, 
    6.592382e-08, 6.612164e-08, 6.410102e-08, 6.422221e-08, 6.421153e-08, 
    6.433836e-08, 6.443215e-08, 6.463544e-08, 6.496149e-08, 6.483888e-08, 
    6.506396e-08, 6.510916e-08, 6.476719e-08, 6.497716e-08, 6.430331e-08, 
    6.441219e-08, 6.434736e-08, 6.411058e-08, 6.486714e-08, 6.447888e-08, 
    6.519582e-08, 6.498549e-08, 6.559934e-08, 6.529407e-08, 6.589367e-08, 
    6.615002e-08, 6.639124e-08, 6.667317e-08, 6.428834e-08, 6.4206e-08, 
    6.435344e-08, 6.455743e-08, 6.47467e-08, 6.499832e-08, 6.502406e-08, 
    6.507121e-08, 6.51933e-08, 6.529596e-08, 6.508611e-08, 6.53217e-08, 
    6.443745e-08, 6.490084e-08, 6.417487e-08, 6.439348e-08, 6.454541e-08, 
    6.447876e-08, 6.482487e-08, 6.490644e-08, 6.523793e-08, 6.506657e-08, 
    6.608675e-08, 6.56354e-08, 6.688783e-08, 6.653783e-08, 6.417723e-08, 
    6.428806e-08, 6.467379e-08, 6.449026e-08, 6.501512e-08, 6.514431e-08, 
    6.524932e-08, 6.538358e-08, 6.539807e-08, 6.547761e-08, 6.534727e-08, 
    6.547247e-08, 6.499886e-08, 6.52105e-08, 6.46297e-08, 6.477106e-08, 
    6.470603e-08, 6.463469e-08, 6.485485e-08, 6.508942e-08, 6.509442e-08, 
    6.516963e-08, 6.53816e-08, 6.501724e-08, 6.614502e-08, 6.544855e-08, 
    6.440892e-08, 6.462241e-08, 6.465289e-08, 6.457019e-08, 6.513136e-08, 
    6.492802e-08, 6.547567e-08, 6.532767e-08, 6.557018e-08, 6.544967e-08, 
    6.543194e-08, 6.527716e-08, 6.51808e-08, 6.493735e-08, 6.473926e-08, 
    6.458218e-08, 6.46187e-08, 6.479126e-08, 6.510376e-08, 6.539939e-08, 
    6.533463e-08, 6.555175e-08, 6.497706e-08, 6.521804e-08, 6.512491e-08, 
    6.536776e-08, 6.483562e-08, 6.528879e-08, 6.471979e-08, 6.476968e-08, 
    6.492399e-08, 6.52344e-08, 6.530306e-08, 6.537638e-08, 6.533113e-08, 
    6.51117e-08, 6.507574e-08, 6.492024e-08, 6.487731e-08, 6.475882e-08, 
    6.466072e-08, 6.475035e-08, 6.484448e-08, 6.511178e-08, 6.535268e-08, 
    6.561532e-08, 6.567959e-08, 6.598647e-08, 6.573666e-08, 6.61489e-08, 
    6.579844e-08, 6.64051e-08, 6.531504e-08, 6.578811e-08, 6.493101e-08, 
    6.502334e-08, 6.519036e-08, 6.557342e-08, 6.536661e-08, 6.560847e-08, 
    6.507433e-08, 6.479721e-08, 6.47255e-08, 6.459173e-08, 6.472857e-08, 
    6.471743e-08, 6.484837e-08, 6.480629e-08, 6.512066e-08, 6.49518e-08, 
    6.54315e-08, 6.560656e-08, 6.610091e-08, 6.640397e-08, 6.671245e-08, 
    6.684864e-08, 6.689009e-08, 6.690742e-08 ;

 LAND_USE_FLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC =
  0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203 ;

 LEAFC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC_LOSS =
  8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10 ;

 LEAFN =
  0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507 ;

 LEAF_MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LFC2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LF_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITFALL =
  1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09 ;

 LITHR =
  8.591897e-13, 8.615078e-13, 8.610575e-13, 8.629254e-13, 8.618897e-13, 
    8.631123e-13, 8.596602e-13, 8.615995e-13, 8.603619e-13, 8.593989e-13, 
    8.66545e-13, 8.630088e-13, 8.702151e-13, 8.679639e-13, 8.736153e-13, 
    8.698645e-13, 8.743711e-13, 8.73508e-13, 8.761065e-13, 8.753624e-13, 
    8.78681e-13, 8.764498e-13, 8.804005e-13, 8.781488e-13, 8.785009e-13, 
    8.76376e-13, 8.637216e-13, 8.661048e-13, 8.635801e-13, 8.639202e-13, 
    8.637678e-13, 8.619109e-13, 8.60974e-13, 8.590129e-13, 8.593692e-13, 
    8.608098e-13, 8.640731e-13, 8.629664e-13, 8.65756e-13, 8.656931e-13, 
    8.687941e-13, 8.673965e-13, 8.726022e-13, 8.711244e-13, 8.753935e-13, 
    8.743204e-13, 8.75343e-13, 8.750331e-13, 8.75347e-13, 8.737731e-13, 
    8.744475e-13, 8.730623e-13, 8.676582e-13, 8.692477e-13, 8.645031e-13, 
    8.616442e-13, 8.597452e-13, 8.58396e-13, 8.585868e-13, 8.589503e-13, 
    8.608182e-13, 8.625737e-13, 8.639103e-13, 8.648039e-13, 8.65684e-13, 
    8.683441e-13, 8.697523e-13, 8.729006e-13, 8.723333e-13, 8.732947e-13, 
    8.742137e-13, 8.757548e-13, 8.755013e-13, 8.761798e-13, 8.732698e-13, 
    8.75204e-13, 8.720105e-13, 8.72884e-13, 8.659207e-13, 8.632651e-13, 
    8.621332e-13, 8.611439e-13, 8.587334e-13, 8.603982e-13, 8.59742e-13, 
    8.613034e-13, 8.622946e-13, 8.618045e-13, 8.648283e-13, 8.636531e-13, 
    8.698358e-13, 8.671749e-13, 8.741065e-13, 8.724498e-13, 8.745035e-13, 
    8.734559e-13, 8.752503e-13, 8.736355e-13, 8.764325e-13, 8.770408e-13, 
    8.766251e-13, 8.782224e-13, 8.735458e-13, 8.753427e-13, 8.617907e-13, 
    8.618706e-13, 8.622432e-13, 8.606048e-13, 8.605048e-13, 8.59003e-13, 
    8.603395e-13, 8.609082e-13, 8.623522e-13, 8.632054e-13, 8.640164e-13, 
    8.657984e-13, 8.677864e-13, 8.70564e-13, 8.725572e-13, 8.738925e-13, 
    8.73074e-13, 8.737966e-13, 8.729887e-13, 8.7261e-13, 8.768127e-13, 
    8.744536e-13, 8.779927e-13, 8.777971e-13, 8.761959e-13, 8.778192e-13, 
    8.619267e-13, 8.614667e-13, 8.598681e-13, 8.611193e-13, 8.588395e-13, 
    8.601155e-13, 8.608488e-13, 8.636771e-13, 8.642987e-13, 8.648741e-13, 
    8.660107e-13, 8.67468e-13, 8.700222e-13, 8.72242e-13, 8.742672e-13, 
    8.74119e-13, 8.741711e-13, 8.746231e-13, 8.735031e-13, 8.748069e-13, 
    8.750254e-13, 8.744537e-13, 8.777709e-13, 8.768238e-13, 8.77793e-13, 
    8.771764e-13, 8.616163e-13, 8.623903e-13, 8.619721e-13, 8.627584e-13, 
    8.622043e-13, 8.646666e-13, 8.654043e-13, 8.688535e-13, 8.674392e-13, 
    8.696903e-13, 8.676682e-13, 8.680265e-13, 8.697626e-13, 8.677777e-13, 
    8.721191e-13, 8.691759e-13, 8.746406e-13, 8.717039e-13, 8.748245e-13, 
    8.742585e-13, 8.751958e-13, 8.760347e-13, 8.7709e-13, 8.79035e-13, 
    8.785849e-13, 8.802109e-13, 8.63544e-13, 8.645469e-13, 8.644591e-13, 
    8.655085e-13, 8.66284e-13, 8.679648e-13, 8.706572e-13, 8.696453e-13, 
    8.715032e-13, 8.718759e-13, 8.690534e-13, 8.707863e-13, 8.652181e-13, 
    8.661182e-13, 8.655827e-13, 8.636229e-13, 8.698778e-13, 8.666697e-13, 
    8.725901e-13, 8.708555e-13, 8.75915e-13, 8.733995e-13, 8.783369e-13, 
    8.804428e-13, 8.824252e-13, 8.847366e-13, 8.650945e-13, 8.644133e-13, 
    8.656333e-13, 8.673193e-13, 8.688838e-13, 8.709612e-13, 8.71174e-13, 
    8.715628e-13, 8.725696e-13, 8.73416e-13, 8.716852e-13, 8.736282e-13, 
    8.663259e-13, 8.701563e-13, 8.641552e-13, 8.659634e-13, 8.672201e-13, 
    8.666694e-13, 8.695298e-13, 8.702032e-13, 8.729369e-13, 8.715247e-13, 
    8.799228e-13, 8.762111e-13, 8.864965e-13, 8.83627e-13, 8.641751e-13, 
    8.650924e-13, 8.682811e-13, 8.667646e-13, 8.711001e-13, 8.721653e-13, 
    8.730316e-13, 8.741377e-13, 8.742575e-13, 8.749126e-13, 8.738389e-13, 
    8.748704e-13, 8.709657e-13, 8.727113e-13, 8.679175e-13, 8.690851e-13, 
    8.685482e-13, 8.679588e-13, 8.697773e-13, 8.717123e-13, 8.717544e-13, 
    8.723739e-13, 8.741185e-13, 8.711177e-13, 8.803999e-13, 8.746705e-13, 
    8.660921e-13, 8.67856e-13, 8.681088e-13, 8.674256e-13, 8.720589e-13, 
    8.703811e-13, 8.748967e-13, 8.736773e-13, 8.756752e-13, 8.746825e-13, 
    8.745364e-13, 8.73261e-13, 8.724663e-13, 8.704579e-13, 8.688223e-13, 
    8.675248e-13, 8.678266e-13, 8.692517e-13, 8.718308e-13, 8.742679e-13, 
    8.737341e-13, 8.755234e-13, 8.70786e-13, 8.727731e-13, 8.720053e-13, 
    8.740076e-13, 8.696182e-13, 8.733541e-13, 8.686619e-13, 8.690739e-13, 
    8.703478e-13, 8.729073e-13, 8.734744e-13, 8.740784e-13, 8.737059e-13, 
    8.718964e-13, 8.716001e-13, 8.703171e-13, 8.699623e-13, 8.689842e-13, 
    8.681739e-13, 8.689141e-13, 8.696911e-13, 8.718975e-13, 8.73883e-13, 
    8.760465e-13, 8.765759e-13, 8.790982e-13, 8.77044e-13, 8.804316e-13, 
    8.775502e-13, 8.825364e-13, 8.735716e-13, 8.77467e-13, 8.70406e-13, 
    8.711681e-13, 8.725444e-13, 8.757007e-13, 8.739981e-13, 8.759895e-13, 
    8.715886e-13, 8.693005e-13, 8.68709e-13, 8.676036e-13, 8.687343e-13, 
    8.686424e-13, 8.697238e-13, 8.693764e-13, 8.719707e-13, 8.705776e-13, 
    8.745325e-13, 8.75974e-13, 8.800403e-13, 8.825286e-13, 8.850598e-13, 
    8.861758e-13, 8.865154e-13, 8.866573e-13 ;

 LITR1C =
  3.066802e-05, 3.066791e-05, 3.066793e-05, 3.066783e-05, 3.066788e-05, 
    3.066782e-05, 3.0668e-05, 3.06679e-05, 3.066796e-05, 3.066801e-05, 
    3.066765e-05, 3.066783e-05, 3.066747e-05, 3.066758e-05, 3.06673e-05, 
    3.066748e-05, 3.066726e-05, 3.06673e-05, 3.066717e-05, 3.066721e-05, 
    3.066704e-05, 3.066715e-05, 3.066696e-05, 3.066707e-05, 3.066705e-05, 
    3.066716e-05, 3.066779e-05, 3.066767e-05, 3.06678e-05, 3.066778e-05, 
    3.066779e-05, 3.066788e-05, 3.066793e-05, 3.066803e-05, 3.066801e-05, 
    3.066794e-05, 3.066778e-05, 3.066783e-05, 3.066769e-05, 3.06677e-05, 
    3.066754e-05, 3.066761e-05, 3.066735e-05, 3.066742e-05, 3.066721e-05, 
    3.066726e-05, 3.066721e-05, 3.066723e-05, 3.066721e-05, 3.066729e-05, 
    3.066726e-05, 3.066732e-05, 3.06676e-05, 3.066752e-05, 3.066775e-05, 
    3.06679e-05, 3.066799e-05, 3.066806e-05, 3.066805e-05, 3.066803e-05, 
    3.066794e-05, 3.066785e-05, 3.066778e-05, 3.066774e-05, 3.06677e-05, 
    3.066756e-05, 3.066749e-05, 3.066733e-05, 3.066736e-05, 3.066731e-05, 
    3.066727e-05, 3.066719e-05, 3.06672e-05, 3.066717e-05, 3.066731e-05, 
    3.066722e-05, 3.066738e-05, 3.066733e-05, 3.066768e-05, 3.066782e-05, 
    3.066787e-05, 3.066792e-05, 3.066804e-05, 3.066796e-05, 3.066799e-05, 
    3.066791e-05, 3.066787e-05, 3.066789e-05, 3.066774e-05, 3.06678e-05, 
    3.066749e-05, 3.066762e-05, 3.066727e-05, 3.066735e-05, 3.066725e-05, 
    3.066731e-05, 3.066722e-05, 3.06673e-05, 3.066715e-05, 3.066712e-05, 
    3.066715e-05, 3.066707e-05, 3.06673e-05, 3.066721e-05, 3.066789e-05, 
    3.066789e-05, 3.066787e-05, 3.066795e-05, 3.066795e-05, 3.066803e-05, 
    3.066796e-05, 3.066794e-05, 3.066786e-05, 3.066782e-05, 3.066778e-05, 
    3.066769e-05, 3.066759e-05, 3.066745e-05, 3.066735e-05, 3.066728e-05, 
    3.066732e-05, 3.066729e-05, 3.066733e-05, 3.066735e-05, 3.066714e-05, 
    3.066726e-05, 3.066708e-05, 3.066709e-05, 3.066717e-05, 3.066708e-05, 
    3.066788e-05, 3.066791e-05, 3.066799e-05, 3.066792e-05, 3.066804e-05, 
    3.066798e-05, 3.066794e-05, 3.06678e-05, 3.066776e-05, 3.066774e-05, 
    3.066768e-05, 3.06676e-05, 3.066748e-05, 3.066736e-05, 3.066726e-05, 
    3.066727e-05, 3.066727e-05, 3.066724e-05, 3.06673e-05, 3.066724e-05, 
    3.066723e-05, 3.066726e-05, 3.066709e-05, 3.066714e-05, 3.066709e-05, 
    3.066712e-05, 3.06679e-05, 3.066786e-05, 3.066788e-05, 3.066784e-05, 
    3.066787e-05, 3.066775e-05, 3.066771e-05, 3.066754e-05, 3.066761e-05, 
    3.06675e-05, 3.066759e-05, 3.066758e-05, 3.066749e-05, 3.066759e-05, 
    3.066737e-05, 3.066752e-05, 3.066724e-05, 3.066739e-05, 3.066724e-05, 
    3.066726e-05, 3.066722e-05, 3.066718e-05, 3.066712e-05, 3.066702e-05, 
    3.066705e-05, 3.066696e-05, 3.06678e-05, 3.066775e-05, 3.066776e-05, 
    3.06677e-05, 3.066767e-05, 3.066758e-05, 3.066744e-05, 3.06675e-05, 
    3.06674e-05, 3.066738e-05, 3.066752e-05, 3.066744e-05, 3.066772e-05, 
    3.066767e-05, 3.06677e-05, 3.06678e-05, 3.066748e-05, 3.066764e-05, 
    3.066735e-05, 3.066743e-05, 3.066718e-05, 3.066731e-05, 3.066706e-05, 
    3.066695e-05, 3.066686e-05, 3.066674e-05, 3.066772e-05, 3.066776e-05, 
    3.06677e-05, 3.066761e-05, 3.066754e-05, 3.066743e-05, 3.066742e-05, 
    3.06674e-05, 3.066735e-05, 3.066731e-05, 3.066739e-05, 3.06673e-05, 
    3.066766e-05, 3.066747e-05, 3.066777e-05, 3.066768e-05, 3.066762e-05, 
    3.066764e-05, 3.06675e-05, 3.066747e-05, 3.066733e-05, 3.06674e-05, 
    3.066698e-05, 3.066716e-05, 3.066665e-05, 3.066679e-05, 3.066777e-05, 
    3.066772e-05, 3.066756e-05, 3.066764e-05, 3.066742e-05, 3.066737e-05, 
    3.066732e-05, 3.066727e-05, 3.066726e-05, 3.066723e-05, 3.066728e-05, 
    3.066723e-05, 3.066743e-05, 3.066734e-05, 3.066758e-05, 3.066752e-05, 
    3.066755e-05, 3.066758e-05, 3.066749e-05, 3.066739e-05, 3.066739e-05, 
    3.066736e-05, 3.066727e-05, 3.066742e-05, 3.066696e-05, 3.066724e-05, 
    3.066767e-05, 3.066759e-05, 3.066757e-05, 3.066761e-05, 3.066738e-05, 
    3.066746e-05, 3.066723e-05, 3.066729e-05, 3.066719e-05, 3.066724e-05, 
    3.066725e-05, 3.066731e-05, 3.066735e-05, 3.066746e-05, 3.066754e-05, 
    3.06676e-05, 3.066759e-05, 3.066752e-05, 3.066739e-05, 3.066726e-05, 
    3.066729e-05, 3.06672e-05, 3.066744e-05, 3.066734e-05, 3.066738e-05, 
    3.066728e-05, 3.06675e-05, 3.066731e-05, 3.066755e-05, 3.066752e-05, 
    3.066746e-05, 3.066733e-05, 3.06673e-05, 3.066727e-05, 3.066729e-05, 
    3.066738e-05, 3.06674e-05, 3.066746e-05, 3.066748e-05, 3.066753e-05, 
    3.066757e-05, 3.066753e-05, 3.06675e-05, 3.066738e-05, 3.066728e-05, 
    3.066718e-05, 3.066715e-05, 3.066702e-05, 3.066712e-05, 3.066695e-05, 
    3.06671e-05, 3.066685e-05, 3.06673e-05, 3.06671e-05, 3.066746e-05, 
    3.066742e-05, 3.066735e-05, 3.066719e-05, 3.066728e-05, 3.066718e-05, 
    3.06674e-05, 3.066751e-05, 3.066754e-05, 3.06676e-05, 3.066754e-05, 
    3.066755e-05, 3.066749e-05, 3.066751e-05, 3.066738e-05, 3.066745e-05, 
    3.066725e-05, 3.066718e-05, 3.066698e-05, 3.066685e-05, 3.066672e-05, 
    3.066667e-05, 3.066665e-05, 3.066664e-05 ;

 LITR1C_TO_SOIL1C =
  5.722613e-13, 5.738049e-13, 5.735051e-13, 5.74749e-13, 5.740592e-13, 
    5.748734e-13, 5.725745e-13, 5.73866e-13, 5.730418e-13, 5.724006e-13, 
    5.771593e-13, 5.748045e-13, 5.796034e-13, 5.781042e-13, 5.818677e-13, 
    5.793699e-13, 5.823709e-13, 5.817962e-13, 5.835266e-13, 5.830311e-13, 
    5.85241e-13, 5.837552e-13, 5.86386e-13, 5.848866e-13, 5.851211e-13, 
    5.837061e-13, 5.752792e-13, 5.768662e-13, 5.75185e-13, 5.754115e-13, 
    5.753099e-13, 5.740733e-13, 5.734495e-13, 5.721435e-13, 5.723808e-13, 
    5.733401e-13, 5.755133e-13, 5.747763e-13, 5.76634e-13, 5.765921e-13, 
    5.786571e-13, 5.777264e-13, 5.81193e-13, 5.802089e-13, 5.830518e-13, 
    5.823372e-13, 5.830181e-13, 5.828117e-13, 5.830208e-13, 5.819727e-13, 
    5.824219e-13, 5.814994e-13, 5.779006e-13, 5.789591e-13, 5.757996e-13, 
    5.738957e-13, 5.726311e-13, 5.717327e-13, 5.718598e-13, 5.721018e-13, 
    5.733457e-13, 5.745147e-13, 5.754048e-13, 5.759999e-13, 5.76586e-13, 
    5.783574e-13, 5.792952e-13, 5.813917e-13, 5.81014e-13, 5.816541e-13, 
    5.822661e-13, 5.832924e-13, 5.831236e-13, 5.835755e-13, 5.816376e-13, 
    5.829256e-13, 5.80799e-13, 5.813806e-13, 5.767436e-13, 5.749752e-13, 
    5.742214e-13, 5.735626e-13, 5.719574e-13, 5.730661e-13, 5.726291e-13, 
    5.736688e-13, 5.743289e-13, 5.740025e-13, 5.760162e-13, 5.752335e-13, 
    5.793508e-13, 5.775788e-13, 5.821948e-13, 5.810915e-13, 5.824591e-13, 
    5.817615e-13, 5.829565e-13, 5.818811e-13, 5.837437e-13, 5.841487e-13, 
    5.838719e-13, 5.849356e-13, 5.818214e-13, 5.83018e-13, 5.739933e-13, 
    5.740465e-13, 5.742946e-13, 5.732036e-13, 5.73137e-13, 5.72137e-13, 
    5.73027e-13, 5.734057e-13, 5.743673e-13, 5.749354e-13, 5.754755e-13, 
    5.766621e-13, 5.77986e-13, 5.798357e-13, 5.81163e-13, 5.820523e-13, 
    5.815072e-13, 5.819884e-13, 5.814504e-13, 5.811982e-13, 5.839969e-13, 
    5.824259e-13, 5.847827e-13, 5.846524e-13, 5.835861e-13, 5.846671e-13, 
    5.740839e-13, 5.737776e-13, 5.72713e-13, 5.735462e-13, 5.72028e-13, 
    5.728778e-13, 5.733661e-13, 5.752495e-13, 5.756635e-13, 5.760466e-13, 
    5.768035e-13, 5.77774e-13, 5.794749e-13, 5.809531e-13, 5.823018e-13, 
    5.822031e-13, 5.822378e-13, 5.825387e-13, 5.817929e-13, 5.826611e-13, 
    5.828066e-13, 5.824259e-13, 5.84635e-13, 5.840043e-13, 5.846497e-13, 
    5.84239e-13, 5.738772e-13, 5.743927e-13, 5.741142e-13, 5.746378e-13, 
    5.742688e-13, 5.759085e-13, 5.763997e-13, 5.786967e-13, 5.777548e-13, 
    5.792539e-13, 5.779073e-13, 5.781459e-13, 5.79302e-13, 5.779802e-13, 
    5.808713e-13, 5.789113e-13, 5.825504e-13, 5.805948e-13, 5.826729e-13, 
    5.822959e-13, 5.829202e-13, 5.834787e-13, 5.841815e-13, 5.854768e-13, 
    5.85177e-13, 5.862598e-13, 5.751609e-13, 5.758287e-13, 5.757703e-13, 
    5.764691e-13, 5.769856e-13, 5.781048e-13, 5.798978e-13, 5.79224e-13, 
    5.804612e-13, 5.807093e-13, 5.788297e-13, 5.799838e-13, 5.762757e-13, 
    5.768751e-13, 5.765185e-13, 5.752134e-13, 5.793788e-13, 5.772424e-13, 
    5.811849e-13, 5.800298e-13, 5.833991e-13, 5.81724e-13, 5.850119e-13, 
    5.864142e-13, 5.877343e-13, 5.892736e-13, 5.761934e-13, 5.757398e-13, 
    5.765523e-13, 5.77675e-13, 5.787168e-13, 5.801003e-13, 5.802419e-13, 
    5.805008e-13, 5.811713e-13, 5.817349e-13, 5.805823e-13, 5.818762e-13, 
    5.770135e-13, 5.795642e-13, 5.755679e-13, 5.76772e-13, 5.776089e-13, 
    5.772422e-13, 5.79147e-13, 5.795955e-13, 5.814159e-13, 5.804754e-13, 
    5.86068e-13, 5.835962e-13, 5.904455e-13, 5.885346e-13, 5.755811e-13, 
    5.76192e-13, 5.783155e-13, 5.773056e-13, 5.801927e-13, 5.80902e-13, 
    5.814789e-13, 5.822155e-13, 5.822953e-13, 5.827316e-13, 5.820165e-13, 
    5.827034e-13, 5.801032e-13, 5.812657e-13, 5.780733e-13, 5.788508e-13, 
    5.784933e-13, 5.781008e-13, 5.793118e-13, 5.806004e-13, 5.806284e-13, 
    5.81041e-13, 5.822027e-13, 5.802044e-13, 5.863856e-13, 5.825703e-13, 
    5.768578e-13, 5.780324e-13, 5.782007e-13, 5.777458e-13, 5.808312e-13, 
    5.79714e-13, 5.82721e-13, 5.819089e-13, 5.832393e-13, 5.825784e-13, 
    5.824811e-13, 5.816317e-13, 5.811025e-13, 5.797651e-13, 5.786759e-13, 
    5.778118e-13, 5.780128e-13, 5.789618e-13, 5.806793e-13, 5.823023e-13, 
    5.819468e-13, 5.831383e-13, 5.799835e-13, 5.813068e-13, 5.807955e-13, 
    5.821289e-13, 5.792059e-13, 5.816937e-13, 5.78569e-13, 5.788434e-13, 
    5.796917e-13, 5.813962e-13, 5.817738e-13, 5.82176e-13, 5.81928e-13, 
    5.80723e-13, 5.805256e-13, 5.796712e-13, 5.79435e-13, 5.787837e-13, 
    5.78244e-13, 5.78737e-13, 5.792544e-13, 5.807237e-13, 5.820459e-13, 
    5.834866e-13, 5.838391e-13, 5.855188e-13, 5.841509e-13, 5.864068e-13, 
    5.84488e-13, 5.878084e-13, 5.818385e-13, 5.844326e-13, 5.797305e-13, 
    5.80238e-13, 5.811545e-13, 5.832564e-13, 5.821226e-13, 5.834487e-13, 
    5.805179e-13, 5.789943e-13, 5.786004e-13, 5.778643e-13, 5.786173e-13, 
    5.78556e-13, 5.792762e-13, 5.790448e-13, 5.807725e-13, 5.798448e-13, 
    5.824785e-13, 5.834384e-13, 5.861462e-13, 5.878032e-13, 5.894888e-13, 
    5.90232e-13, 5.904581e-13, 5.905526e-13 ;

 LITR1C_vr =
  0.001751176, 0.001751169, 0.00175117, 0.001751165, 0.001751168, 
    0.001751164, 0.001751174, 0.001751169, 0.001751172, 0.001751175, 
    0.001751155, 0.001751165, 0.001751144, 0.001751151, 0.001751134, 
    0.001751145, 0.001751132, 0.001751135, 0.001751127, 0.001751129, 
    0.00175112, 0.001751126, 0.001751115, 0.001751121, 0.00175112, 
    0.001751126, 0.001751163, 0.001751156, 0.001751163, 0.001751162, 
    0.001751163, 0.001751168, 0.001751171, 0.001751176, 0.001751175, 
    0.001751171, 0.001751162, 0.001751165, 0.001751157, 0.001751157, 
    0.001751148, 0.001751152, 0.001751137, 0.001751142, 0.001751129, 
    0.001751132, 0.001751129, 0.00175113, 0.001751129, 0.001751134, 
    0.001751132, 0.001751136, 0.001751151, 0.001751147, 0.00175116, 
    0.001751169, 0.001751174, 0.001751178, 0.001751177, 0.001751176, 
    0.001751171, 0.001751166, 0.001751162, 0.00175116, 0.001751157, 
    0.001751149, 0.001751145, 0.001751136, 0.001751138, 0.001751135, 
    0.001751133, 0.001751128, 0.001751129, 0.001751127, 0.001751135, 
    0.00175113, 0.001751139, 0.001751136, 0.001751156, 0.001751164, 
    0.001751167, 0.00175117, 0.001751177, 0.001751172, 0.001751174, 
    0.00175117, 0.001751167, 0.001751168, 0.00175116, 0.001751163, 
    0.001751145, 0.001751153, 0.001751133, 0.001751138, 0.001751132, 
    0.001751135, 0.00175113, 0.001751134, 0.001751126, 0.001751125, 
    0.001751126, 0.001751121, 0.001751135, 0.001751129, 0.001751168, 
    0.001751168, 0.001751167, 0.001751172, 0.001751172, 0.001751176, 
    0.001751172, 0.001751171, 0.001751167, 0.001751164, 0.001751162, 
    0.001751157, 0.001751151, 0.001751143, 0.001751137, 0.001751134, 
    0.001751136, 0.001751134, 0.001751136, 0.001751137, 0.001751125, 
    0.001751132, 0.001751122, 0.001751122, 0.001751127, 0.001751122, 
    0.001751168, 0.001751169, 0.001751174, 0.00175117, 0.001751177, 
    0.001751173, 0.001751171, 0.001751163, 0.001751161, 0.001751159, 
    0.001751156, 0.001751152, 0.001751145, 0.001751138, 0.001751132, 
    0.001751133, 0.001751133, 0.001751131, 0.001751135, 0.001751131, 
    0.00175113, 0.001751132, 0.001751122, 0.001751125, 0.001751122, 
    0.001751124, 0.001751169, 0.001751167, 0.001751168, 0.001751165, 
    0.001751167, 0.00175116, 0.001751158, 0.001751148, 0.001751152, 
    0.001751146, 0.001751151, 0.00175115, 0.001751145, 0.001751151, 
    0.001751139, 0.001751147, 0.001751131, 0.00175114, 0.001751131, 
    0.001751133, 0.00175113, 0.001751127, 0.001751124, 0.001751119, 
    0.00175112, 0.001751115, 0.001751163, 0.00175116, 0.001751161, 
    0.001751158, 0.001751155, 0.001751151, 0.001751143, 0.001751146, 
    0.00175114, 0.001751139, 0.001751147, 0.001751142, 0.001751158, 
    0.001751156, 0.001751157, 0.001751163, 0.001751145, 0.001751154, 
    0.001751137, 0.001751142, 0.001751128, 0.001751135, 0.001751121, 
    0.001751115, 0.001751109, 0.001751102, 0.001751159, 0.001751161, 
    0.001751157, 0.001751152, 0.001751148, 0.001751142, 0.001751141, 
    0.00175114, 0.001751137, 0.001751135, 0.00175114, 0.001751134, 
    0.001751155, 0.001751144, 0.001751162, 0.001751156, 0.001751153, 
    0.001751154, 0.001751146, 0.001751144, 0.001751136, 0.00175114, 
    0.001751116, 0.001751127, 0.001751097, 0.001751106, 0.001751161, 
    0.001751159, 0.00175115, 0.001751154, 0.001751142, 0.001751138, 
    0.001751136, 0.001751133, 0.001751133, 0.001751131, 0.001751134, 
    0.001751131, 0.001751142, 0.001751137, 0.001751151, 0.001751147, 
    0.001751149, 0.001751151, 0.001751145, 0.00175114, 0.00175114, 
    0.001751138, 0.001751133, 0.001751142, 0.001751115, 0.001751131, 
    0.001751156, 0.001751151, 0.00175115, 0.001751152, 0.001751139, 
    0.001751144, 0.001751131, 0.001751134, 0.001751128, 0.001751131, 
    0.001751132, 0.001751135, 0.001751138, 0.001751143, 0.001751148, 
    0.001751152, 0.001751151, 0.001751147, 0.001751139, 0.001751132, 
    0.001751134, 0.001751129, 0.001751142, 0.001751137, 0.001751139, 
    0.001751133, 0.001751146, 0.001751135, 0.001751148, 0.001751147, 
    0.001751144, 0.001751136, 0.001751135, 0.001751133, 0.001751134, 
    0.001751139, 0.00175114, 0.001751144, 0.001751145, 0.001751148, 
    0.00175115, 0.001751148, 0.001751146, 0.001751139, 0.001751134, 
    0.001751127, 0.001751126, 0.001751119, 0.001751125, 0.001751115, 
    0.001751123, 0.001751109, 0.001751134, 0.001751123, 0.001751143, 
    0.001751141, 0.001751137, 0.001751128, 0.001751133, 0.001751128, 
    0.00175114, 0.001751147, 0.001751148, 0.001751152, 0.001751148, 
    0.001751149, 0.001751145, 0.001751147, 0.001751139, 0.001751143, 
    0.001751132, 0.001751128, 0.001751116, 0.001751109, 0.001751101, 
    0.001751098, 0.001751097, 0.001751097,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N =
  9.73289e-07, 9.732854e-07, 9.732861e-07, 9.732831e-07, 9.732847e-07, 
    9.732828e-07, 9.732884e-07, 9.732853e-07, 9.732872e-07, 9.732887e-07, 
    9.732773e-07, 9.73283e-07, 9.732715e-07, 9.732751e-07, 9.732661e-07, 
    9.732721e-07, 9.732648e-07, 9.732663e-07, 9.732621e-07, 9.732632e-07, 
    9.73258e-07, 9.732615e-07, 9.732553e-07, 9.732588e-07, 9.732582e-07, 
    9.732616e-07, 9.732819e-07, 9.73278e-07, 9.732821e-07, 9.732815e-07, 
    9.732818e-07, 9.732847e-07, 9.732862e-07, 9.732894e-07, 9.732888e-07, 
    9.732865e-07, 9.732813e-07, 9.73283e-07, 9.732786e-07, 9.732787e-07, 
    9.732738e-07, 9.73276e-07, 9.732677e-07, 9.732701e-07, 9.732632e-07, 
    9.732649e-07, 9.732634e-07, 9.732638e-07, 9.732634e-07, 9.732659e-07, 
    9.732647e-07, 9.73267e-07, 9.732756e-07, 9.73273e-07, 9.732806e-07, 
    9.732852e-07, 9.732883e-07, 9.732904e-07, 9.732901e-07, 9.732895e-07, 
    9.732865e-07, 9.732837e-07, 9.732815e-07, 9.732802e-07, 9.732787e-07, 
    9.732745e-07, 9.732722e-07, 9.732672e-07, 9.732681e-07, 9.732665e-07, 
    9.732652e-07, 9.732627e-07, 9.732631e-07, 9.73262e-07, 9.732667e-07, 
    9.732636e-07, 9.732687e-07, 9.732672e-07, 9.732784e-07, 9.732826e-07, 
    9.732844e-07, 9.73286e-07, 9.732898e-07, 9.732871e-07, 9.732883e-07, 
    9.732858e-07, 9.732842e-07, 9.73285e-07, 9.732801e-07, 9.73282e-07, 
    9.732721e-07, 9.732763e-07, 9.732653e-07, 9.732679e-07, 9.732647e-07, 
    9.732663e-07, 9.732635e-07, 9.732661e-07, 9.732615e-07, 9.732606e-07, 
    9.732613e-07, 9.732587e-07, 9.732662e-07, 9.732634e-07, 9.73285e-07, 
    9.732848e-07, 9.732843e-07, 9.732869e-07, 9.73287e-07, 9.732894e-07, 
    9.732872e-07, 9.732863e-07, 9.73284e-07, 9.732827e-07, 9.732814e-07, 
    9.732786e-07, 9.732754e-07, 9.73271e-07, 9.732678e-07, 9.732656e-07, 
    9.73267e-07, 9.732657e-07, 9.732671e-07, 9.732677e-07, 9.73261e-07, 
    9.732647e-07, 9.732591e-07, 9.732594e-07, 9.73262e-07, 9.732594e-07, 
    9.732847e-07, 9.732854e-07, 9.73288e-07, 9.73286e-07, 9.732896e-07, 
    9.732876e-07, 9.732864e-07, 9.732819e-07, 9.73281e-07, 9.732801e-07, 
    9.732782e-07, 9.732759e-07, 9.732718e-07, 9.732682e-07, 9.732651e-07, 
    9.732653e-07, 9.732652e-07, 9.732645e-07, 9.732663e-07, 9.732642e-07, 
    9.732638e-07, 9.732647e-07, 9.732595e-07, 9.73261e-07, 9.732594e-07, 
    9.732604e-07, 9.732852e-07, 9.732839e-07, 9.732846e-07, 9.732834e-07, 
    9.732843e-07, 9.732804e-07, 9.732792e-07, 9.732737e-07, 9.73276e-07, 
    9.732723e-07, 9.732755e-07, 9.73275e-07, 9.732722e-07, 9.732754e-07, 
    9.732685e-07, 9.732731e-07, 9.732645e-07, 9.732692e-07, 9.732642e-07, 
    9.732651e-07, 9.732636e-07, 9.732622e-07, 9.732605e-07, 9.732574e-07, 
    9.732581e-07, 9.732556e-07, 9.732821e-07, 9.732805e-07, 9.732806e-07, 
    9.73279e-07, 9.732778e-07, 9.732751e-07, 9.732707e-07, 9.732724e-07, 
    9.732695e-07, 9.732688e-07, 9.732734e-07, 9.732706e-07, 9.732795e-07, 
    9.73278e-07, 9.732789e-07, 9.73282e-07, 9.73272e-07, 9.732771e-07, 
    9.732677e-07, 9.732705e-07, 9.732624e-07, 9.732664e-07, 9.732586e-07, 
    9.732552e-07, 9.73252e-07, 9.732483e-07, 9.732797e-07, 9.732807e-07, 
    9.732788e-07, 9.732761e-07, 9.732736e-07, 9.732703e-07, 9.732699e-07, 
    9.732694e-07, 9.732678e-07, 9.732664e-07, 9.732692e-07, 9.732661e-07, 
    9.732777e-07, 9.732717e-07, 9.732812e-07, 9.732782e-07, 9.732763e-07, 
    9.732771e-07, 9.732726e-07, 9.732715e-07, 9.732672e-07, 9.732694e-07, 
    9.732561e-07, 9.73262e-07, 9.732455e-07, 9.732502e-07, 9.732811e-07, 
    9.732797e-07, 9.732746e-07, 9.73277e-07, 9.732701e-07, 9.732684e-07, 
    9.73267e-07, 9.732653e-07, 9.732651e-07, 9.73264e-07, 9.732657e-07, 
    9.73264e-07, 9.732703e-07, 9.732676e-07, 9.732752e-07, 9.732734e-07, 
    9.732742e-07, 9.732751e-07, 9.732722e-07, 9.732692e-07, 9.73269e-07, 
    9.73268e-07, 9.732653e-07, 9.732701e-07, 9.732553e-07, 9.732644e-07, 
    9.732781e-07, 9.732753e-07, 9.732748e-07, 9.73276e-07, 9.732686e-07, 
    9.732712e-07, 9.73264e-07, 9.73266e-07, 9.732628e-07, 9.732644e-07, 
    9.732646e-07, 9.732667e-07, 9.732679e-07, 9.732711e-07, 9.732737e-07, 
    9.732757e-07, 9.732753e-07, 9.73273e-07, 9.732689e-07, 9.732651e-07, 
    9.732659e-07, 9.73263e-07, 9.732706e-07, 9.732674e-07, 9.732687e-07, 
    9.732654e-07, 9.732724e-07, 9.732665e-07, 9.732739e-07, 9.732734e-07, 
    9.732713e-07, 9.732672e-07, 9.732663e-07, 9.732653e-07, 9.73266e-07, 
    9.732688e-07, 9.732693e-07, 9.732713e-07, 9.732719e-07, 9.732735e-07, 
    9.732747e-07, 9.732736e-07, 9.732723e-07, 9.732688e-07, 9.732656e-07, 
    9.732622e-07, 9.732613e-07, 9.732573e-07, 9.732606e-07, 9.732552e-07, 
    9.732598e-07, 9.732519e-07, 9.732662e-07, 9.732599e-07, 9.732712e-07, 
    9.732699e-07, 9.732678e-07, 9.732628e-07, 9.732655e-07, 9.732623e-07, 
    9.732693e-07, 9.73273e-07, 9.732739e-07, 9.732756e-07, 9.732738e-07, 
    9.73274e-07, 9.732723e-07, 9.732728e-07, 9.732687e-07, 9.73271e-07, 
    9.732646e-07, 9.732623e-07, 9.732559e-07, 9.732519e-07, 9.732479e-07, 
    9.732461e-07, 9.732455e-07, 9.732453e-07 ;

 LITR1N_TNDNCY_VERT_TRANS =
  1.470543e-25, 4.362612e-25, -1.960724e-26, 3.333231e-25, -3.725376e-25, 
    1.078398e-25, -2.156797e-25, -4.019485e-25, -1.323489e-25, 3.333231e-25, 
    6.862535e-26, -9.313441e-26, 1.240158e-24, -4.901811e-26, 9.019333e-25, 
    -1.274471e-25, 2.205815e-25, -3.039123e-25, 7.646825e-25, 2.548942e-25, 
    5.931191e-25, -4.41163e-26, 5.342974e-25, -7.352717e-26, 2.548942e-25, 
    -3.823413e-25, 4.362612e-25, -6.078246e-25, -1.960724e-26, -2.646978e-25, 
    5.391992e-25, -3.333231e-25, 1.666616e-25, -1.068595e-24, 3.872431e-25, 
    -9.803622e-26, 8.82326e-26, 7.548789e-25, -1.960724e-26, -4.901811e-26, 
    2.548942e-25, 3.823413e-25, -3.921449e-25, 2.941087e-25, 1.421525e-25, 
    2.843051e-25, 3.039123e-25, -5.686101e-25, -7.842898e-26, -2.450906e-25, 
    2.548942e-25, 4.313593e-25, -5.588064e-25, 4.65672e-25, 5.19592e-25, 
    4.019485e-25, 4.558684e-25, -1.56858e-25, -5.882173e-25, 8.235043e-25, 
    -1.127417e-25, -4.999847e-25, 6.421373e-25, -3.529304e-25, -5.784137e-25, 
    -1.960724e-26, 3.480286e-25, 1.323489e-25, -4.509666e-25, -7.842898e-26, 
    9.803622e-27, 1.24506e-24, 5.833155e-25, 4.019485e-25, 2.843051e-25, 
    8.725224e-25, -3.137159e-25, 5.882173e-25, 3.333231e-25, 3.039123e-25, 
    -3.088141e-25, -1.960724e-25, 2.646978e-25, 4.117521e-25, -1.470543e-25, 
    5.98021e-25, 0, 6.078246e-25, -4.803775e-25, -4.901811e-25, 3.235195e-25, 
    1.02938e-25, 1.176435e-25, -2.156797e-25, 2.352869e-25, -1.421525e-25, 
    6.862535e-26, -3.529304e-25, -3.137159e-25, 3.137159e-25, 9.999695e-25, 
    9.803622e-26, 0, 5.490028e-25, 6.421373e-25, 3.333231e-25, 4.264576e-25, 
    -5.882173e-25, 3.529304e-25, 4.019485e-25, -2.499924e-25, -1.56858e-25, 
    -3.039123e-25, 6.862535e-25, 1.127417e-25, -1.372507e-24, 9.313441e-25, 
    -3.62734e-25, 7.352717e-26, 4.313593e-25, -9.999695e-25, -3.725376e-25, 
    -6.421373e-25, 6.372354e-26, 2.303851e-25, 3.823413e-25, 6.960572e-25, 
    -3.431268e-25, -5.097883e-25, 1.088202e-24, -6.274318e-25, -3.186177e-25, 
    -4.65672e-25, -5.490028e-25, -1.470543e-25, 8.921296e-25, 7.646825e-25, 
    9.803622e-26, 3.774394e-25, -6.176282e-25, 2.59796e-25, -7.058608e-25, 
    -5.882173e-26, 9.803622e-26, 2.695996e-25, 2.156797e-25, -8.137007e-25, 
    4.950829e-25, -6.862535e-26, 6.372354e-25, -2.058761e-25, 3.725376e-25, 
    5.490028e-25, 2.058761e-25, 6.568427e-25, 1.862688e-25, 3.088141e-25, 
    3.431268e-25, 7.79388e-25, 1.470543e-25, 4.901811e-25, 3.137159e-25, 
    2.254833e-25, 2.450905e-26, -2.401887e-25, -4.607703e-25, 4.901811e-25, 
    4.754757e-25, 7.25468e-25, -1.960724e-26, -9.019333e-25, 5.588064e-25, 
    2.352869e-25, 3.529304e-25, 1.960724e-25, -9.313441e-26, -6.122413e-41, 
    -1.274471e-25, -3.137159e-25, 8.725224e-25, 4.901811e-26, -4.705739e-25, 
    -6.47039e-25, -4.803775e-25, 3.62734e-25, 2.352869e-25, 6.372354e-25, 
    6.2253e-25, -1.470543e-25, 1.176435e-25, -2.009742e-25, -4.117521e-25, 
    -1.960724e-26, 3.235195e-25, -4.803775e-25, 3.186177e-25, 2.352869e-25, 
    7.058608e-25, 3.529304e-25, 2.450906e-25, 6.568427e-25, -5.048866e-25, 
    1.372507e-25, -6.862535e-26, -4.607703e-25, -1.372507e-25, -1.862688e-25, 
    -7.450753e-25, 1.004871e-24, -4.068503e-25, -9.60755e-25, -8.333079e-26, 
    -1.372507e-25, -3.431268e-25, 4.705739e-25, -2.254833e-25, 6.813517e-25, 
    -3.676358e-25, 3.137159e-25, 8.725224e-25, -4.068503e-25, -6.122413e-41, 
    -2.941087e-26, 7.352717e-26, 2.205815e-25, 4.754757e-25, 8.137007e-25, 
    5.686101e-25, 6.274318e-25, 2.058761e-25, 8.627187e-25, 2.156797e-25, 
    6.47039e-25, 4.019485e-25, -5.882173e-26, 1.274471e-25, -3.431268e-25, 
    -1.323489e-25, 2.450905e-26, 2.843051e-25, -2.450906e-25, 4.313593e-25, 
    6.274318e-25, -9.803622e-26, -6.274318e-25, 9.803622e-26, -2.401887e-25, 
    8.82326e-26, 2.548942e-25, 5.391992e-26, 4.509666e-25, 5.882173e-25, 
    -1.56858e-25, 1.078398e-25, 8.235043e-25, 9.215405e-25, 0, -3.235195e-25, 
    -3.725376e-25, -9.803622e-26, 3.529304e-25, 1.004871e-24, 2.450905e-26, 
    -5.490028e-25, -6.078246e-25, 5.097883e-25, 6.862535e-26, -5.931191e-25, 
    2.59796e-25, 3.137159e-25, 8.82326e-26, 1.421525e-25, 6.519409e-25, 
    -3.431268e-26, -7.107626e-25, 9.803622e-27, -9.803622e-25, -2.548942e-25, 
    -6.372354e-26, 2.058761e-25, 3.333231e-25, 5.490028e-25, -6.274318e-25, 
    2.058761e-25, -4.901811e-25, 9.117368e-25, -6.862535e-26, 3.235195e-25, 
    -2.941087e-25, 7.156644e-25, -4.117521e-25, 4.264576e-25, -6.47039e-25, 
    -9.509513e-25, 5.19592e-25, 4.215557e-25, -1.156827e-24, 2.303851e-25, 
    1.470543e-25, -1.862688e-25, 6.176282e-25, -4.117521e-25, 5.686101e-25, 
    3.970467e-25, 1.911706e-25, -1.960724e-26, 4.901811e-26, 2.254833e-25, 
    -1.960724e-25, -1.519561e-25, -4.901811e-26, 3.921449e-25, 9.803622e-26, 
    -3.431268e-25, 5.735119e-25, -2.548942e-25, -2.352869e-25, 1.127417e-25, 
    7.352717e-25, 4.215557e-25, -4.705739e-25, 3.039123e-25, 9.803622e-26, 
    2.941087e-26, -6.274318e-25, 1.666616e-25, -3.872431e-25, 7.352717e-25, 
    7.25468e-25, -2.352869e-25, -3.529304e-25, -4.901811e-26, 5.391992e-26, 
    -6.078246e-25, 8.82326e-26, 3.039123e-25, 2.745014e-25, -2.254833e-25,
  9.436731e-32, 9.436693e-32, 9.436701e-32, 9.436671e-32, 9.436688e-32, 
    9.436668e-32, 9.436723e-32, 9.436692e-32, 9.436712e-32, 9.436728e-32, 
    9.436613e-32, 9.436669e-32, 9.436554e-32, 9.43659e-32, 9.4365e-32, 
    9.436559e-32, 9.436487e-32, 9.436501e-32, 9.43646e-32, 9.436471e-32, 
    9.436418e-32, 9.436454e-32, 9.436391e-32, 9.436427e-32, 9.436421e-32, 
    9.436455e-32, 9.436658e-32, 9.43662e-32, 9.436661e-32, 9.436655e-32, 
    9.436658e-32, 9.436687e-32, 9.436702e-32, 9.436733e-32, 9.436728e-32, 
    9.436705e-32, 9.436652e-32, 9.43667e-32, 9.436625e-32, 9.436626e-32, 
    9.436577e-32, 9.436599e-32, 9.436516e-32, 9.43654e-32, 9.436471e-32, 
    9.436488e-32, 9.436472e-32, 9.436477e-32, 9.436472e-32, 9.436497e-32, 
    9.436486e-32, 9.436508e-32, 9.436595e-32, 9.436569e-32, 9.436645e-32, 
    9.436691e-32, 9.436722e-32, 9.436743e-32, 9.436741e-32, 9.436735e-32, 
    9.436705e-32, 9.436676e-32, 9.436655e-32, 9.436641e-32, 9.436626e-32, 
    9.436584e-32, 9.436561e-32, 9.436511e-32, 9.43652e-32, 9.436505e-32, 
    9.43649e-32, 9.436465e-32, 9.43647e-32, 9.436458e-32, 9.436505e-32, 
    9.436474e-32, 9.436525e-32, 9.436511e-32, 9.436623e-32, 9.436665e-32, 
    9.436684e-32, 9.436699e-32, 9.436738e-32, 9.436711e-32, 9.436722e-32, 
    9.436697e-32, 9.436681e-32, 9.436689e-32, 9.436641e-32, 9.436659e-32, 
    9.43656e-32, 9.436603e-32, 9.436492e-32, 9.436518e-32, 9.436485e-32, 
    9.436502e-32, 9.436473e-32, 9.4365e-32, 9.436454e-32, 9.436445e-32, 
    9.436451e-32, 9.436426e-32, 9.436501e-32, 9.436472e-32, 9.436689e-32, 
    9.436688e-32, 9.436682e-32, 9.436708e-32, 9.436709e-32, 9.436733e-32, 
    9.436712e-32, 9.436703e-32, 9.43668e-32, 9.436666e-32, 9.436654e-32, 
    9.436625e-32, 9.436593e-32, 9.436548e-32, 9.436517e-32, 9.436495e-32, 
    9.436508e-32, 9.436497e-32, 9.43651e-32, 9.436515e-32, 9.436448e-32, 
    9.436486e-32, 9.43643e-32, 9.436433e-32, 9.436458e-32, 9.436433e-32, 
    9.436687e-32, 9.436694e-32, 9.43672e-32, 9.4367e-32, 9.436736e-32, 
    9.436716e-32, 9.436704e-32, 9.436659e-32, 9.436649e-32, 9.436639e-32, 
    9.436621e-32, 9.436598e-32, 9.436557e-32, 9.436521e-32, 9.436489e-32, 
    9.436491e-32, 9.436491e-32, 9.436484e-32, 9.436501e-32, 9.436481e-32, 
    9.436477e-32, 9.436486e-32, 9.436433e-32, 9.436448e-32, 9.436433e-32, 
    9.436443e-32, 9.436692e-32, 9.436679e-32, 9.436686e-32, 9.436674e-32, 
    9.436682e-32, 9.436643e-32, 9.436631e-32, 9.436576e-32, 9.436598e-32, 
    9.436562e-32, 9.436595e-32, 9.436589e-32, 9.436561e-32, 9.436593e-32, 
    9.436524e-32, 9.436571e-32, 9.436483e-32, 9.43653e-32, 9.43648e-32, 
    9.43649e-32, 9.436474e-32, 9.436461e-32, 9.436444e-32, 9.436413e-32, 
    9.43642e-32, 9.436394e-32, 9.436661e-32, 9.436645e-32, 9.436646e-32, 
    9.436629e-32, 9.436617e-32, 9.43659e-32, 9.436547e-32, 9.436563e-32, 
    9.436534e-32, 9.436527e-32, 9.436572e-32, 9.436545e-32, 9.436634e-32, 
    9.436619e-32, 9.436628e-32, 9.436659e-32, 9.436559e-32, 9.436611e-32, 
    9.436516e-32, 9.436544e-32, 9.436463e-32, 9.436503e-32, 9.436424e-32, 
    9.43639e-32, 9.436358e-32, 9.436321e-32, 9.436636e-32, 9.436647e-32, 
    9.436628e-32, 9.436601e-32, 9.436575e-32, 9.436542e-32, 9.436539e-32, 
    9.436532e-32, 9.436517e-32, 9.436502e-32, 9.436531e-32, 9.4365e-32, 
    9.436617e-32, 9.436555e-32, 9.436651e-32, 9.436622e-32, 9.436602e-32, 
    9.436611e-32, 9.436565e-32, 9.436554e-32, 9.436511e-32, 9.436533e-32, 
    9.436398e-32, 9.436458e-32, 9.436293e-32, 9.436339e-32, 9.436651e-32, 
    9.436636e-32, 9.436585e-32, 9.436609e-32, 9.43654e-32, 9.436523e-32, 
    9.436509e-32, 9.436491e-32, 9.43649e-32, 9.436479e-32, 9.436496e-32, 
    9.43648e-32, 9.436542e-32, 9.436514e-32, 9.436591e-32, 9.436572e-32, 
    9.436581e-32, 9.43659e-32, 9.436561e-32, 9.43653e-32, 9.43653e-32, 
    9.43652e-32, 9.436491e-32, 9.43654e-32, 9.436391e-32, 9.436482e-32, 
    9.43662e-32, 9.436592e-32, 9.436588e-32, 9.436599e-32, 9.436524e-32, 
    9.436551e-32, 9.436479e-32, 9.436498e-32, 9.436467e-32, 9.436482e-32, 
    9.436485e-32, 9.436505e-32, 9.436518e-32, 9.43655e-32, 9.436577e-32, 
    9.436597e-32, 9.436592e-32, 9.436569e-32, 9.436528e-32, 9.436489e-32, 
    9.436498e-32, 9.436469e-32, 9.436545e-32, 9.436513e-32, 9.436525e-32, 
    9.436493e-32, 9.436564e-32, 9.436504e-32, 9.436579e-32, 9.436572e-32, 
    9.436552e-32, 9.436511e-32, 9.436502e-32, 9.436492e-32, 9.436498e-32, 
    9.436527e-32, 9.436532e-32, 9.436552e-32, 9.436558e-32, 9.436574e-32, 
    9.436587e-32, 9.436575e-32, 9.436562e-32, 9.436527e-32, 9.436495e-32, 
    9.436461e-32, 9.436452e-32, 9.436412e-32, 9.436445e-32, 9.43639e-32, 
    9.436437e-32, 9.436357e-32, 9.4365e-32, 9.436438e-32, 9.436551e-32, 
    9.436539e-32, 9.436517e-32, 9.436466e-32, 9.436494e-32, 9.436461e-32, 
    9.436532e-32, 9.436569e-32, 9.436578e-32, 9.436596e-32, 9.436578e-32, 
    9.436579e-32, 9.436562e-32, 9.436568e-32, 9.436526e-32, 9.436548e-32, 
    9.436485e-32, 9.436462e-32, 9.436397e-32, 9.436357e-32, 9.436316e-32, 
    9.436299e-32, 9.436293e-32, 9.436291e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N_TO_SOIL1N =
  4.035863e-14, 4.04675e-14, 4.044635e-14, 4.053407e-14, 4.048543e-14, 
    4.054285e-14, 4.038072e-14, 4.04718e-14, 4.041368e-14, 4.036846e-14, 
    4.070406e-14, 4.053799e-14, 4.087643e-14, 4.07707e-14, 4.103612e-14, 
    4.085996e-14, 4.107161e-14, 4.103108e-14, 4.115312e-14, 4.111817e-14, 
    4.127402e-14, 4.116924e-14, 4.135478e-14, 4.124903e-14, 4.126556e-14, 
    4.116577e-14, 4.057147e-14, 4.068339e-14, 4.056482e-14, 4.05808e-14, 
    4.057364e-14, 4.048643e-14, 4.044243e-14, 4.035033e-14, 4.036706e-14, 
    4.043472e-14, 4.058798e-14, 4.0536e-14, 4.066701e-14, 4.066406e-14, 
    4.08097e-14, 4.074406e-14, 4.098854e-14, 4.091914e-14, 4.111963e-14, 
    4.106923e-14, 4.111726e-14, 4.11027e-14, 4.111745e-14, 4.104353e-14, 
    4.10752e-14, 4.101014e-14, 4.075635e-14, 4.0831e-14, 4.060817e-14, 
    4.04739e-14, 4.038471e-14, 4.032135e-14, 4.033032e-14, 4.034738e-14, 
    4.043511e-14, 4.051756e-14, 4.058033e-14, 4.062229e-14, 4.066363e-14, 
    4.078856e-14, 4.08547e-14, 4.100255e-14, 4.097591e-14, 4.102106e-14, 
    4.106422e-14, 4.11366e-14, 4.112469e-14, 4.115656e-14, 4.101989e-14, 
    4.111073e-14, 4.096075e-14, 4.100177e-14, 4.067475e-14, 4.055003e-14, 
    4.049687e-14, 4.045041e-14, 4.03372e-14, 4.041539e-14, 4.038457e-14, 
    4.04579e-14, 4.050445e-14, 4.048143e-14, 4.062344e-14, 4.056825e-14, 
    4.085862e-14, 4.073365e-14, 4.105919e-14, 4.098138e-14, 4.107783e-14, 
    4.102863e-14, 4.111291e-14, 4.103707e-14, 4.116843e-14, 4.119699e-14, 
    4.117747e-14, 4.125249e-14, 4.103285e-14, 4.111725e-14, 4.048078e-14, 
    4.048454e-14, 4.050203e-14, 4.042509e-14, 4.042039e-14, 4.034986e-14, 
    4.041263e-14, 4.043934e-14, 4.050716e-14, 4.054723e-14, 4.058531e-14, 
    4.0669e-14, 4.076237e-14, 4.089282e-14, 4.098643e-14, 4.104914e-14, 
    4.10107e-14, 4.104463e-14, 4.100669e-14, 4.098891e-14, 4.118628e-14, 
    4.107549e-14, 4.12417e-14, 4.123251e-14, 4.115731e-14, 4.123355e-14, 
    4.048717e-14, 4.046557e-14, 4.039049e-14, 4.044925e-14, 4.034218e-14, 
    4.040211e-14, 4.043655e-14, 4.056938e-14, 4.059857e-14, 4.062559e-14, 
    4.067897e-14, 4.074742e-14, 4.086737e-14, 4.097162e-14, 4.106674e-14, 
    4.105977e-14, 4.106222e-14, 4.108345e-14, 4.103085e-14, 4.109208e-14, 
    4.110234e-14, 4.107549e-14, 4.123128e-14, 4.11868e-14, 4.123232e-14, 
    4.120336e-14, 4.047259e-14, 4.050895e-14, 4.04893e-14, 4.052623e-14, 
    4.050021e-14, 4.061585e-14, 4.065049e-14, 4.081248e-14, 4.074606e-14, 
    4.085179e-14, 4.075682e-14, 4.077364e-14, 4.085518e-14, 4.076196e-14, 
    4.096585e-14, 4.082763e-14, 4.108427e-14, 4.094635e-14, 4.109291e-14, 
    4.106633e-14, 4.111034e-14, 4.114974e-14, 4.11993e-14, 4.129065e-14, 
    4.126951e-14, 4.134588e-14, 4.056313e-14, 4.061023e-14, 4.06061e-14, 
    4.065539e-14, 4.069181e-14, 4.077075e-14, 4.08972e-14, 4.084967e-14, 
    4.093693e-14, 4.095443e-14, 4.082187e-14, 4.090325e-14, 4.064175e-14, 
    4.068402e-14, 4.065887e-14, 4.056683e-14, 4.086059e-14, 4.070992e-14, 
    4.098797e-14, 4.09065e-14, 4.114412e-14, 4.102598e-14, 4.125786e-14, 
    4.135677e-14, 4.144987e-14, 4.155842e-14, 4.063594e-14, 4.060395e-14, 
    4.066125e-14, 4.074043e-14, 4.081391e-14, 4.091147e-14, 4.092146e-14, 
    4.093972e-14, 4.098701e-14, 4.102676e-14, 4.094547e-14, 4.103672e-14, 
    4.069378e-14, 4.087367e-14, 4.059183e-14, 4.067675e-14, 4.073577e-14, 
    4.070991e-14, 4.084424e-14, 4.087587e-14, 4.100426e-14, 4.093794e-14, 
    4.133234e-14, 4.115803e-14, 4.164107e-14, 4.150631e-14, 4.059276e-14, 
    4.063585e-14, 4.07856e-14, 4.071438e-14, 4.091799e-14, 4.096802e-14, 
    4.10087e-14, 4.106065e-14, 4.106628e-14, 4.109705e-14, 4.104662e-14, 
    4.109506e-14, 4.091168e-14, 4.099366e-14, 4.076852e-14, 4.082336e-14, 
    4.079814e-14, 4.077046e-14, 4.085587e-14, 4.094674e-14, 4.094872e-14, 
    4.097782e-14, 4.105975e-14, 4.091882e-14, 4.135475e-14, 4.108568e-14, 
    4.06828e-14, 4.076564e-14, 4.077751e-14, 4.074542e-14, 4.096302e-14, 
    4.088423e-14, 4.10963e-14, 4.103903e-14, 4.113286e-14, 4.108624e-14, 
    4.107938e-14, 4.101948e-14, 4.098216e-14, 4.088784e-14, 4.081102e-14, 
    4.075008e-14, 4.076426e-14, 4.083118e-14, 4.095231e-14, 4.106677e-14, 
    4.10417e-14, 4.112573e-14, 4.090324e-14, 4.099656e-14, 4.096051e-14, 
    4.105454e-14, 4.08484e-14, 4.102385e-14, 4.080348e-14, 4.082283e-14, 
    4.088266e-14, 4.100287e-14, 4.10295e-14, 4.105787e-14, 4.104037e-14, 
    4.095539e-14, 4.094147e-14, 4.088122e-14, 4.086456e-14, 4.081863e-14, 
    4.078056e-14, 4.081533e-14, 4.085182e-14, 4.095544e-14, 4.104869e-14, 
    4.11503e-14, 4.117516e-14, 4.129362e-14, 4.119714e-14, 4.135624e-14, 
    4.122092e-14, 4.145509e-14, 4.103406e-14, 4.121701e-14, 4.08854e-14, 
    4.092119e-14, 4.098583e-14, 4.113405e-14, 4.10541e-14, 4.114762e-14, 
    4.094093e-14, 4.083347e-14, 4.08057e-14, 4.075378e-14, 4.080689e-14, 
    4.080257e-14, 4.085336e-14, 4.083704e-14, 4.095888e-14, 4.089345e-14, 
    4.10792e-14, 4.114689e-14, 4.133786e-14, 4.145472e-14, 4.15736e-14, 
    4.162601e-14, 4.164196e-14, 4.164863e-14 ;

 LITR1N_vr =
  5.557581e-05, 5.55756e-05, 5.557564e-05, 5.557547e-05, 5.557557e-05, 
    5.557546e-05, 5.557577e-05, 5.557559e-05, 5.557571e-05, 5.557579e-05, 
    5.557514e-05, 5.557546e-05, 5.557481e-05, 5.557501e-05, 5.55745e-05, 
    5.557484e-05, 5.557443e-05, 5.557451e-05, 5.557427e-05, 5.557434e-05, 
    5.557404e-05, 5.557424e-05, 5.557388e-05, 5.557409e-05, 5.557406e-05, 
    5.557425e-05, 5.55754e-05, 5.557518e-05, 5.557541e-05, 5.557538e-05, 
    5.557539e-05, 5.557557e-05, 5.557565e-05, 5.557583e-05, 5.55758e-05, 
    5.557567e-05, 5.557537e-05, 5.557547e-05, 5.557522e-05, 5.557522e-05, 
    5.557494e-05, 5.557507e-05, 5.557459e-05, 5.557472e-05, 5.557434e-05, 
    5.557443e-05, 5.557434e-05, 5.557437e-05, 5.557434e-05, 5.557448e-05, 
    5.557442e-05, 5.557455e-05, 5.557504e-05, 5.55749e-05, 5.557533e-05, 
    5.557559e-05, 5.557576e-05, 5.557589e-05, 5.557587e-05, 5.557583e-05, 
    5.557566e-05, 5.55755e-05, 5.557538e-05, 5.55753e-05, 5.557522e-05, 
    5.557498e-05, 5.557485e-05, 5.557456e-05, 5.557462e-05, 5.557453e-05, 
    5.557444e-05, 5.55743e-05, 5.557433e-05, 5.557427e-05, 5.557453e-05, 
    5.557435e-05, 5.557464e-05, 5.557456e-05, 5.55752e-05, 5.557544e-05, 
    5.557554e-05, 5.557563e-05, 5.557586e-05, 5.55757e-05, 5.557576e-05, 
    5.557562e-05, 5.557553e-05, 5.557558e-05, 5.55753e-05, 5.55754e-05, 
    5.557484e-05, 5.557508e-05, 5.557446e-05, 5.55746e-05, 5.557442e-05, 
    5.557451e-05, 5.557435e-05, 5.55745e-05, 5.557424e-05, 5.557419e-05, 
    5.557423e-05, 5.557408e-05, 5.557451e-05, 5.557434e-05, 5.557558e-05, 
    5.557557e-05, 5.557554e-05, 5.557569e-05, 5.557569e-05, 5.557583e-05, 
    5.557571e-05, 5.557566e-05, 5.557553e-05, 5.557545e-05, 5.557537e-05, 
    5.557521e-05, 5.557503e-05, 5.557478e-05, 5.557459e-05, 5.557447e-05, 
    5.557455e-05, 5.557448e-05, 5.557456e-05, 5.557459e-05, 5.557421e-05, 
    5.557442e-05, 5.55741e-05, 5.557412e-05, 5.557426e-05, 5.557412e-05, 
    5.557557e-05, 5.557561e-05, 5.557575e-05, 5.557564e-05, 5.557585e-05, 
    5.557573e-05, 5.557566e-05, 5.55754e-05, 5.557535e-05, 5.55753e-05, 
    5.557519e-05, 5.557506e-05, 5.557483e-05, 5.557462e-05, 5.557444e-05, 
    5.557445e-05, 5.557445e-05, 5.557441e-05, 5.557451e-05, 5.557439e-05, 
    5.557437e-05, 5.557442e-05, 5.557412e-05, 5.557421e-05, 5.557412e-05, 
    5.557418e-05, 5.557559e-05, 5.557552e-05, 5.557556e-05, 5.557549e-05, 
    5.557554e-05, 5.557531e-05, 5.557524e-05, 5.557493e-05, 5.557506e-05, 
    5.557486e-05, 5.557504e-05, 5.557501e-05, 5.557485e-05, 5.557503e-05, 
    5.557463e-05, 5.55749e-05, 5.55744e-05, 5.557467e-05, 5.557439e-05, 
    5.557444e-05, 5.557435e-05, 5.557428e-05, 5.557418e-05, 5.5574e-05, 
    5.557405e-05, 5.55739e-05, 5.557542e-05, 5.557532e-05, 5.557533e-05, 
    5.557524e-05, 5.557516e-05, 5.557501e-05, 5.557477e-05, 5.557486e-05, 
    5.557469e-05, 5.557466e-05, 5.557491e-05, 5.557476e-05, 5.557526e-05, 
    5.557518e-05, 5.557523e-05, 5.557541e-05, 5.557484e-05, 5.557513e-05, 
    5.557459e-05, 5.557475e-05, 5.557429e-05, 5.557452e-05, 5.557407e-05, 
    5.557388e-05, 5.55737e-05, 5.557349e-05, 5.557527e-05, 5.557534e-05, 
    5.557523e-05, 5.557507e-05, 5.557493e-05, 5.557474e-05, 5.557472e-05, 
    5.557468e-05, 5.557459e-05, 5.557452e-05, 5.557467e-05, 5.55745e-05, 
    5.557516e-05, 5.557482e-05, 5.557536e-05, 5.557519e-05, 5.557508e-05, 
    5.557513e-05, 5.557487e-05, 5.557481e-05, 5.557456e-05, 5.557469e-05, 
    5.557392e-05, 5.557426e-05, 5.557333e-05, 5.557359e-05, 5.557536e-05, 
    5.557527e-05, 5.557498e-05, 5.557512e-05, 5.557473e-05, 5.557463e-05, 
    5.557455e-05, 5.557445e-05, 5.557444e-05, 5.557438e-05, 5.557448e-05, 
    5.557439e-05, 5.557474e-05, 5.557458e-05, 5.557502e-05, 5.557491e-05, 
    5.557496e-05, 5.557502e-05, 5.557485e-05, 5.557467e-05, 5.557467e-05, 
    5.557461e-05, 5.557445e-05, 5.557472e-05, 5.557388e-05, 5.55744e-05, 
    5.557518e-05, 5.557502e-05, 5.5575e-05, 5.557506e-05, 5.557464e-05, 
    5.557479e-05, 5.557438e-05, 5.557449e-05, 5.557431e-05, 5.55744e-05, 
    5.557442e-05, 5.557453e-05, 5.55746e-05, 5.557479e-05, 5.557494e-05, 
    5.557505e-05, 5.557503e-05, 5.55749e-05, 5.557466e-05, 5.557444e-05, 
    5.557449e-05, 5.557432e-05, 5.557476e-05, 5.557458e-05, 5.557464e-05, 
    5.557446e-05, 5.557486e-05, 5.557452e-05, 5.557495e-05, 5.557491e-05, 
    5.55748e-05, 5.557456e-05, 5.557451e-05, 5.557446e-05, 5.557449e-05, 
    5.557466e-05, 5.557468e-05, 5.55748e-05, 5.557483e-05, 5.557492e-05, 
    5.557499e-05, 5.557493e-05, 5.557486e-05, 5.557466e-05, 5.557447e-05, 
    5.557428e-05, 5.557423e-05, 5.5574e-05, 5.557419e-05, 5.557388e-05, 
    5.557414e-05, 5.557369e-05, 5.55745e-05, 5.557415e-05, 5.557479e-05, 
    5.557472e-05, 5.55746e-05, 5.557431e-05, 5.557446e-05, 5.557428e-05, 
    5.557468e-05, 5.557489e-05, 5.557495e-05, 5.557504e-05, 5.557494e-05, 
    5.557495e-05, 5.557485e-05, 5.557488e-05, 5.557465e-05, 5.557478e-05, 
    5.557442e-05, 5.557428e-05, 5.557391e-05, 5.557369e-05, 5.557346e-05, 
    5.557336e-05, 5.557332e-05, 5.557331e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1_HR =
  6.994304e-13, 7.013172e-13, 7.009506e-13, 7.02471e-13, 7.01628e-13, 
    7.026231e-13, 6.998134e-13, 7.013917e-13, 7.003845e-13, 6.996007e-13, 
    7.05417e-13, 7.025388e-13, 7.084041e-13, 7.065718e-13, 7.111716e-13, 
    7.081188e-13, 7.117866e-13, 7.110842e-13, 7.131991e-13, 7.125936e-13, 
    7.152945e-13, 7.134786e-13, 7.166941e-13, 7.148614e-13, 7.15148e-13, 
    7.134185e-13, 7.03119e-13, 7.050587e-13, 7.030038e-13, 7.032806e-13, 
    7.031566e-13, 7.016452e-13, 7.008827e-13, 6.992865e-13, 6.995765e-13, 
    7.00749e-13, 7.034051e-13, 7.025043e-13, 7.047749e-13, 7.047237e-13, 
    7.072476e-13, 7.0611e-13, 7.10347e-13, 7.091442e-13, 7.126189e-13, 
    7.117455e-13, 7.125777e-13, 7.123255e-13, 7.12581e-13, 7.112999e-13, 
    7.118489e-13, 7.107214e-13, 7.06323e-13, 7.076167e-13, 7.037551e-13, 
    7.014282e-13, 6.998825e-13, 6.987845e-13, 6.989397e-13, 6.992355e-13, 
    7.007559e-13, 7.021847e-13, 7.032726e-13, 7.039998e-13, 7.047162e-13, 
    7.068813e-13, 7.080275e-13, 7.105898e-13, 7.101281e-13, 7.109106e-13, 
    7.116586e-13, 7.129129e-13, 7.127066e-13, 7.132589e-13, 7.108904e-13, 
    7.124646e-13, 7.098654e-13, 7.105763e-13, 7.049089e-13, 7.027475e-13, 
    7.018262e-13, 7.01021e-13, 6.99059e-13, 7.004141e-13, 6.9988e-13, 
    7.011508e-13, 7.019575e-13, 7.015587e-13, 7.040197e-13, 7.030633e-13, 
    7.080954e-13, 7.059297e-13, 7.115714e-13, 7.10223e-13, 7.118945e-13, 
    7.110418e-13, 7.125024e-13, 7.11188e-13, 7.134645e-13, 7.139596e-13, 
    7.136212e-13, 7.149213e-13, 7.11115e-13, 7.125775e-13, 7.015474e-13, 
    7.016124e-13, 7.019157e-13, 7.005822e-13, 7.005007e-13, 6.992785e-13, 
    7.003663e-13, 7.008292e-13, 7.020044e-13, 7.026989e-13, 7.033589e-13, 
    7.048093e-13, 7.064273e-13, 7.08688e-13, 7.103104e-13, 7.113972e-13, 
    7.10731e-13, 7.113191e-13, 7.106616e-13, 7.103534e-13, 7.13774e-13, 
    7.118539e-13, 7.147344e-13, 7.145752e-13, 7.132719e-13, 7.145932e-13, 
    7.016581e-13, 7.012837e-13, 6.999826e-13, 7.010009e-13, 6.991454e-13, 
    7.00184e-13, 7.007807e-13, 7.030828e-13, 7.035887e-13, 7.04057e-13, 
    7.049821e-13, 7.061683e-13, 7.082471e-13, 7.100538e-13, 7.117022e-13, 
    7.115815e-13, 7.11624e-13, 7.119918e-13, 7.110802e-13, 7.121414e-13, 
    7.123193e-13, 7.118539e-13, 7.145539e-13, 7.13783e-13, 7.145718e-13, 
    7.1407e-13, 7.014055e-13, 7.020355e-13, 7.01695e-13, 7.023351e-13, 
    7.01884e-13, 7.038881e-13, 7.044885e-13, 7.072959e-13, 7.061448e-13, 
    7.07977e-13, 7.063312e-13, 7.066228e-13, 7.080358e-13, 7.064203e-13, 
    7.099538e-13, 7.075583e-13, 7.120061e-13, 7.096158e-13, 7.121558e-13, 
    7.116951e-13, 7.124579e-13, 7.131407e-13, 7.139996e-13, 7.155827e-13, 
    7.152164e-13, 7.165398e-13, 7.029745e-13, 7.037907e-13, 7.037192e-13, 
    7.045733e-13, 7.052046e-13, 7.065726e-13, 7.08764e-13, 7.079404e-13, 
    7.094526e-13, 7.097558e-13, 7.074586e-13, 7.08869e-13, 7.04337e-13, 
    7.050696e-13, 7.046338e-13, 7.030386e-13, 7.081296e-13, 7.055185e-13, 
    7.103371e-13, 7.089253e-13, 7.130433e-13, 7.109959e-13, 7.150145e-13, 
    7.167285e-13, 7.183419e-13, 7.202233e-13, 7.042364e-13, 7.03682e-13, 
    7.04675e-13, 7.060472e-13, 7.073205e-13, 7.090114e-13, 7.091846e-13, 
    7.09501e-13, 7.103205e-13, 7.110093e-13, 7.096006e-13, 7.11182e-13, 
    7.052387e-13, 7.083563e-13, 7.034719e-13, 7.049436e-13, 7.059665e-13, 
    7.055183e-13, 7.078463e-13, 7.083944e-13, 7.106194e-13, 7.0947e-13, 
    7.163053e-13, 7.132842e-13, 7.216556e-13, 7.193201e-13, 7.034881e-13, 
    7.042347e-13, 7.0683e-13, 7.055957e-13, 7.091244e-13, 7.099914e-13, 
    7.106965e-13, 7.115967e-13, 7.116942e-13, 7.122274e-13, 7.113536e-13, 
    7.121931e-13, 7.09015e-13, 7.104358e-13, 7.065341e-13, 7.074844e-13, 
    7.070474e-13, 7.065677e-13, 7.080478e-13, 7.096227e-13, 7.09657e-13, 
    7.101612e-13, 7.115811e-13, 7.091387e-13, 7.166936e-13, 7.120304e-13, 
    7.050484e-13, 7.06484e-13, 7.066898e-13, 7.061337e-13, 7.099048e-13, 
    7.085392e-13, 7.122146e-13, 7.11222e-13, 7.128481e-13, 7.120402e-13, 
    7.119213e-13, 7.108832e-13, 7.102364e-13, 7.086017e-13, 7.072705e-13, 
    7.062144e-13, 7.064601e-13, 7.0762e-13, 7.097192e-13, 7.117028e-13, 
    7.112683e-13, 7.127246e-13, 7.088688e-13, 7.104861e-13, 7.098612e-13, 
    7.114908e-13, 7.079183e-13, 7.10959e-13, 7.0714e-13, 7.074753e-13, 
    7.085121e-13, 7.105953e-13, 7.110569e-13, 7.115484e-13, 7.112453e-13, 
    7.097725e-13, 7.095313e-13, 7.084871e-13, 7.081984e-13, 7.074023e-13, 
    7.067427e-13, 7.073452e-13, 7.079776e-13, 7.097734e-13, 7.113894e-13, 
    7.131503e-13, 7.135812e-13, 7.156341e-13, 7.139623e-13, 7.167194e-13, 
    7.143742e-13, 7.184325e-13, 7.11136e-13, 7.143065e-13, 7.085595e-13, 
    7.091798e-13, 7.103e-13, 7.128689e-13, 7.114832e-13, 7.131039e-13, 
    7.09522e-13, 7.076597e-13, 7.071783e-13, 7.062786e-13, 7.071989e-13, 
    7.071241e-13, 7.080042e-13, 7.077215e-13, 7.09833e-13, 7.086992e-13, 
    7.119182e-13, 7.130913e-13, 7.164009e-13, 7.184262e-13, 7.204863e-13, 
    7.213946e-13, 7.21671e-13, 7.217866e-13 ;

 LITR2C =
  1.9396e-05, 1.939598e-05, 1.939598e-05, 1.939597e-05, 1.939597e-05, 
    1.939596e-05, 1.939599e-05, 1.939598e-05, 1.939599e-05, 1.939599e-05, 
    1.939593e-05, 1.939597e-05, 1.939591e-05, 1.939592e-05, 1.939588e-05, 
    1.939591e-05, 1.939587e-05, 1.939588e-05, 1.939585e-05, 1.939586e-05, 
    1.939583e-05, 1.939585e-05, 1.939582e-05, 1.939584e-05, 1.939583e-05, 
    1.939585e-05, 1.939596e-05, 1.939594e-05, 1.939596e-05, 1.939596e-05, 
    1.939596e-05, 1.939597e-05, 1.939598e-05, 1.9396e-05, 1.9396e-05, 
    1.939598e-05, 1.939596e-05, 1.939597e-05, 1.939594e-05, 1.939594e-05, 
    1.939592e-05, 1.939593e-05, 1.939588e-05, 1.93959e-05, 1.939586e-05, 
    1.939587e-05, 1.939586e-05, 1.939586e-05, 1.939586e-05, 1.939587e-05, 
    1.939587e-05, 1.939588e-05, 1.939593e-05, 1.939591e-05, 1.939595e-05, 
    1.939598e-05, 1.939599e-05, 1.9396e-05, 1.9396e-05, 1.9396e-05, 
    1.939598e-05, 1.939597e-05, 1.939596e-05, 1.939595e-05, 1.939594e-05, 
    1.939592e-05, 1.939591e-05, 1.939588e-05, 1.939589e-05, 1.939588e-05, 
    1.939587e-05, 1.939586e-05, 1.939586e-05, 1.939585e-05, 1.939588e-05, 
    1.939586e-05, 1.939589e-05, 1.939588e-05, 1.939594e-05, 1.939596e-05, 
    1.939597e-05, 1.939598e-05, 1.9396e-05, 1.939599e-05, 1.939599e-05, 
    1.939598e-05, 1.939597e-05, 1.939597e-05, 1.939595e-05, 1.939596e-05, 
    1.939591e-05, 1.939593e-05, 1.939587e-05, 1.939589e-05, 1.939587e-05, 
    1.939588e-05, 1.939586e-05, 1.939588e-05, 1.939585e-05, 1.939585e-05, 
    1.939585e-05, 1.939584e-05, 1.939588e-05, 1.939586e-05, 1.939597e-05, 
    1.939597e-05, 1.939597e-05, 1.939599e-05, 1.939599e-05, 1.9396e-05, 
    1.939599e-05, 1.939598e-05, 1.939597e-05, 1.939596e-05, 1.939596e-05, 
    1.939594e-05, 1.939593e-05, 1.93959e-05, 1.939589e-05, 1.939587e-05, 
    1.939588e-05, 1.939587e-05, 1.939588e-05, 1.939588e-05, 1.939585e-05, 
    1.939587e-05, 1.939584e-05, 1.939584e-05, 1.939585e-05, 1.939584e-05, 
    1.939597e-05, 1.939598e-05, 1.939599e-05, 1.939598e-05, 1.9396e-05, 
    1.939599e-05, 1.939598e-05, 1.939596e-05, 1.939595e-05, 1.939595e-05, 
    1.939594e-05, 1.939593e-05, 1.939591e-05, 1.939589e-05, 1.939587e-05, 
    1.939587e-05, 1.939587e-05, 1.939587e-05, 1.939588e-05, 1.939587e-05, 
    1.939586e-05, 1.939587e-05, 1.939584e-05, 1.939585e-05, 1.939584e-05, 
    1.939585e-05, 1.939598e-05, 1.939597e-05, 1.939597e-05, 1.939597e-05, 
    1.939597e-05, 1.939595e-05, 1.939595e-05, 1.939592e-05, 1.939593e-05, 
    1.939591e-05, 1.939593e-05, 1.939592e-05, 1.939591e-05, 1.939593e-05, 
    1.939589e-05, 1.939591e-05, 1.939587e-05, 1.939589e-05, 1.939587e-05, 
    1.939587e-05, 1.939586e-05, 1.939586e-05, 1.939585e-05, 1.939583e-05, 
    1.939583e-05, 1.939582e-05, 1.939596e-05, 1.939595e-05, 1.939595e-05, 
    1.939594e-05, 1.939594e-05, 1.939592e-05, 1.93959e-05, 1.939591e-05, 
    1.939589e-05, 1.939589e-05, 1.939591e-05, 1.93959e-05, 1.939595e-05, 
    1.939594e-05, 1.939594e-05, 1.939596e-05, 1.939591e-05, 1.939593e-05, 
    1.939589e-05, 1.93959e-05, 1.939586e-05, 1.939588e-05, 1.939584e-05, 
    1.939582e-05, 1.93958e-05, 1.939578e-05, 1.939595e-05, 1.939595e-05, 
    1.939594e-05, 1.939593e-05, 1.939592e-05, 1.93959e-05, 1.93959e-05, 
    1.939589e-05, 1.939589e-05, 1.939588e-05, 1.939589e-05, 1.939588e-05, 
    1.939594e-05, 1.939591e-05, 1.939596e-05, 1.939594e-05, 1.939593e-05, 
    1.939593e-05, 1.939591e-05, 1.939591e-05, 1.939588e-05, 1.939589e-05, 
    1.939582e-05, 1.939585e-05, 1.939577e-05, 1.939579e-05, 1.939595e-05, 
    1.939595e-05, 1.939592e-05, 1.939593e-05, 1.93959e-05, 1.939589e-05, 
    1.939588e-05, 1.939587e-05, 1.939587e-05, 1.939587e-05, 1.939587e-05, 
    1.939587e-05, 1.93959e-05, 1.939588e-05, 1.939592e-05, 1.939591e-05, 
    1.939592e-05, 1.939592e-05, 1.939591e-05, 1.939589e-05, 1.939589e-05, 
    1.939589e-05, 1.939587e-05, 1.93959e-05, 1.939582e-05, 1.939587e-05, 
    1.939594e-05, 1.939592e-05, 1.939592e-05, 1.939593e-05, 1.939589e-05, 
    1.93959e-05, 1.939587e-05, 1.939588e-05, 1.939586e-05, 1.939587e-05, 
    1.939587e-05, 1.939588e-05, 1.939589e-05, 1.93959e-05, 1.939592e-05, 
    1.939593e-05, 1.939593e-05, 1.939591e-05, 1.939589e-05, 1.939587e-05, 
    1.939587e-05, 1.939586e-05, 1.93959e-05, 1.939588e-05, 1.939589e-05, 
    1.939587e-05, 1.939591e-05, 1.939588e-05, 1.939592e-05, 1.939591e-05, 
    1.93959e-05, 1.939588e-05, 1.939588e-05, 1.939587e-05, 1.939587e-05, 
    1.939589e-05, 1.939589e-05, 1.93959e-05, 1.939591e-05, 1.939591e-05, 
    1.939592e-05, 1.939592e-05, 1.939591e-05, 1.939589e-05, 1.939587e-05, 
    1.939586e-05, 1.939585e-05, 1.939583e-05, 1.939585e-05, 1.939582e-05, 
    1.939584e-05, 1.93958e-05, 1.939588e-05, 1.939584e-05, 1.93959e-05, 
    1.93959e-05, 1.939589e-05, 1.939586e-05, 1.939587e-05, 1.939586e-05, 
    1.939589e-05, 1.939591e-05, 1.939592e-05, 1.939593e-05, 1.939592e-05, 
    1.939592e-05, 1.939591e-05, 1.939591e-05, 1.939589e-05, 1.93959e-05, 
    1.939587e-05, 1.939586e-05, 1.939582e-05, 1.93958e-05, 1.939578e-05, 
    1.939577e-05, 1.939577e-05, 1.939577e-05 ;

 LITR2C_TO_SOIL1C =
  1.065062e-13, 1.067938e-13, 1.067379e-13, 1.069696e-13, 1.068412e-13, 
    1.069928e-13, 1.065646e-13, 1.068051e-13, 1.066516e-13, 1.065321e-13, 
    1.074187e-13, 1.0698e-13, 1.07874e-13, 1.075947e-13, 1.082958e-13, 
    1.078305e-13, 1.083896e-13, 1.082825e-13, 1.086049e-13, 1.085126e-13, 
    1.089243e-13, 1.086475e-13, 1.091376e-13, 1.088583e-13, 1.089019e-13, 
    1.086383e-13, 1.070684e-13, 1.073641e-13, 1.070509e-13, 1.070931e-13, 
    1.070741e-13, 1.068438e-13, 1.067275e-13, 1.064843e-13, 1.065285e-13, 
    1.067072e-13, 1.07112e-13, 1.069747e-13, 1.073208e-13, 1.07313e-13, 
    1.076977e-13, 1.075243e-13, 1.081701e-13, 1.079868e-13, 1.085164e-13, 
    1.083833e-13, 1.085102e-13, 1.084717e-13, 1.085107e-13, 1.083154e-13, 
    1.083991e-13, 1.082272e-13, 1.075568e-13, 1.07754e-13, 1.071654e-13, 
    1.068107e-13, 1.065751e-13, 1.064077e-13, 1.064314e-13, 1.064765e-13, 
    1.067082e-13, 1.06926e-13, 1.070918e-13, 1.072027e-13, 1.073119e-13, 
    1.076419e-13, 1.078166e-13, 1.082072e-13, 1.081368e-13, 1.082561e-13, 
    1.083701e-13, 1.085613e-13, 1.085298e-13, 1.08614e-13, 1.08253e-13, 
    1.084929e-13, 1.080967e-13, 1.082051e-13, 1.073412e-13, 1.070118e-13, 
    1.068714e-13, 1.067486e-13, 1.064496e-13, 1.066561e-13, 1.065747e-13, 
    1.067684e-13, 1.068914e-13, 1.068306e-13, 1.072057e-13, 1.070599e-13, 
    1.078269e-13, 1.074968e-13, 1.083568e-13, 1.081512e-13, 1.08406e-13, 
    1.082761e-13, 1.084987e-13, 1.082983e-13, 1.086453e-13, 1.087208e-13, 
    1.086692e-13, 1.088674e-13, 1.082872e-13, 1.085101e-13, 1.068289e-13, 
    1.068388e-13, 1.06885e-13, 1.066818e-13, 1.066693e-13, 1.06483e-13, 
    1.066488e-13, 1.067194e-13, 1.068985e-13, 1.070044e-13, 1.07105e-13, 
    1.073261e-13, 1.075727e-13, 1.079173e-13, 1.081646e-13, 1.083302e-13, 
    1.082287e-13, 1.083183e-13, 1.082181e-13, 1.081711e-13, 1.086925e-13, 
    1.083998e-13, 1.088389e-13, 1.088146e-13, 1.08616e-13, 1.088174e-13, 
    1.068457e-13, 1.067887e-13, 1.065903e-13, 1.067456e-13, 1.064627e-13, 
    1.066211e-13, 1.06712e-13, 1.070629e-13, 1.0714e-13, 1.072114e-13, 
    1.073524e-13, 1.075332e-13, 1.078501e-13, 1.081255e-13, 1.083767e-13, 
    1.083583e-13, 1.083648e-13, 1.084209e-13, 1.082819e-13, 1.084437e-13, 
    1.084708e-13, 1.083998e-13, 1.088114e-13, 1.086939e-13, 1.088141e-13, 
    1.087376e-13, 1.068072e-13, 1.069033e-13, 1.068514e-13, 1.069489e-13, 
    1.068802e-13, 1.071856e-13, 1.072772e-13, 1.077051e-13, 1.075296e-13, 
    1.078089e-13, 1.07558e-13, 1.076025e-13, 1.078179e-13, 1.075716e-13, 
    1.081102e-13, 1.077451e-13, 1.08423e-13, 1.080587e-13, 1.084459e-13, 
    1.083756e-13, 1.084919e-13, 1.08596e-13, 1.087269e-13, 1.089682e-13, 
    1.089124e-13, 1.091141e-13, 1.070464e-13, 1.071708e-13, 1.071599e-13, 
    1.072901e-13, 1.073863e-13, 1.075948e-13, 1.079289e-13, 1.078033e-13, 
    1.080338e-13, 1.0808e-13, 1.077299e-13, 1.079449e-13, 1.072541e-13, 
    1.073657e-13, 1.072993e-13, 1.070562e-13, 1.078322e-13, 1.074342e-13, 
    1.081686e-13, 1.079534e-13, 1.085811e-13, 1.082691e-13, 1.088816e-13, 
    1.091429e-13, 1.093888e-13, 1.096756e-13, 1.072387e-13, 1.071542e-13, 
    1.073056e-13, 1.075147e-13, 1.077088e-13, 1.079666e-13, 1.07993e-13, 
    1.080412e-13, 1.081661e-13, 1.082711e-13, 1.080564e-13, 1.082974e-13, 
    1.073915e-13, 1.078667e-13, 1.071222e-13, 1.073465e-13, 1.075024e-13, 
    1.074341e-13, 1.07789e-13, 1.078725e-13, 1.082117e-13, 1.080365e-13, 
    1.090784e-13, 1.086179e-13, 1.098939e-13, 1.095379e-13, 1.071247e-13, 
    1.072385e-13, 1.076341e-13, 1.074459e-13, 1.079838e-13, 1.081159e-13, 
    1.082234e-13, 1.083606e-13, 1.083755e-13, 1.084568e-13, 1.083236e-13, 
    1.084515e-13, 1.079671e-13, 1.081837e-13, 1.07589e-13, 1.077338e-13, 
    1.076672e-13, 1.075941e-13, 1.078197e-13, 1.080597e-13, 1.08065e-13, 
    1.081418e-13, 1.083583e-13, 1.07986e-13, 1.091376e-13, 1.084267e-13, 
    1.073625e-13, 1.075813e-13, 1.076127e-13, 1.075279e-13, 1.081027e-13, 
    1.078946e-13, 1.084548e-13, 1.083035e-13, 1.085514e-13, 1.084282e-13, 
    1.084101e-13, 1.082519e-13, 1.081533e-13, 1.079041e-13, 1.077012e-13, 
    1.075402e-13, 1.075777e-13, 1.077545e-13, 1.080744e-13, 1.083768e-13, 
    1.083106e-13, 1.085326e-13, 1.079448e-13, 1.081913e-13, 1.080961e-13, 
    1.083445e-13, 1.078e-13, 1.082634e-13, 1.076813e-13, 1.077324e-13, 
    1.078905e-13, 1.08208e-13, 1.082784e-13, 1.083533e-13, 1.083071e-13, 
    1.080826e-13, 1.080458e-13, 1.078866e-13, 1.078426e-13, 1.077213e-13, 
    1.076208e-13, 1.077126e-13, 1.07809e-13, 1.080827e-13, 1.08329e-13, 
    1.085975e-13, 1.086631e-13, 1.089761e-13, 1.087212e-13, 1.091415e-13, 
    1.08784e-13, 1.094026e-13, 1.082904e-13, 1.087737e-13, 1.078977e-13, 
    1.079922e-13, 1.08163e-13, 1.085545e-13, 1.083433e-13, 1.085904e-13, 
    1.080444e-13, 1.077605e-13, 1.076872e-13, 1.0755e-13, 1.076903e-13, 
    1.076789e-13, 1.078131e-13, 1.0777e-13, 1.080918e-13, 1.07919e-13, 
    1.084096e-13, 1.085885e-13, 1.090929e-13, 1.094016e-13, 1.097157e-13, 
    1.098541e-13, 1.098963e-13, 1.099139e-13 ;

 LITR2C_vr =
  0.001107531, 0.00110753, 0.001107531, 0.00110753, 0.00110753, 0.00110753, 
    0.001107531, 0.00110753, 0.001107531, 0.001107531, 0.001107528, 
    0.00110753, 0.001107526, 0.001107527, 0.001107525, 0.001107526, 
    0.001107524, 0.001107525, 0.001107523, 0.001107524, 0.001107522, 
    0.001107523, 0.001107521, 0.001107522, 0.001107522, 0.001107523, 
    0.001107529, 0.001107528, 0.001107529, 0.001107529, 0.001107529, 
    0.00110753, 0.001107531, 0.001107532, 0.001107531, 0.001107531, 
    0.001107529, 0.00110753, 0.001107528, 0.001107528, 0.001107527, 
    0.001107528, 0.001107525, 0.001107526, 0.001107524, 0.001107524, 
    0.001107524, 0.001107524, 0.001107524, 0.001107524, 0.001107524, 
    0.001107525, 0.001107527, 0.001107527, 0.001107529, 0.00110753, 
    0.001107531, 0.001107532, 0.001107532, 0.001107532, 0.001107531, 
    0.00110753, 0.001107529, 0.001107529, 0.001107528, 0.001107527, 
    0.001107526, 0.001107525, 0.001107525, 0.001107525, 0.001107524, 
    0.001107524, 0.001107524, 0.001107523, 0.001107525, 0.001107524, 
    0.001107525, 0.001107525, 0.001107528, 0.00110753, 0.00110753, 
    0.001107531, 0.001107532, 0.001107531, 0.001107531, 0.00110753, 
    0.00110753, 0.00110753, 0.001107529, 0.001107529, 0.001107526, 
    0.001107528, 0.001107524, 0.001107525, 0.001107524, 0.001107525, 
    0.001107524, 0.001107525, 0.001107523, 0.001107523, 0.001107523, 
    0.001107522, 0.001107525, 0.001107524, 0.00110753, 0.00110753, 
    0.00110753, 0.001107531, 0.001107531, 0.001107532, 0.001107531, 
    0.001107531, 0.00110753, 0.00110753, 0.001107529, 0.001107528, 
    0.001107527, 0.001107526, 0.001107525, 0.001107524, 0.001107525, 
    0.001107524, 0.001107525, 0.001107525, 0.001107523, 0.001107524, 
    0.001107523, 0.001107523, 0.001107523, 0.001107523, 0.00110753, 
    0.00110753, 0.001107531, 0.001107531, 0.001107532, 0.001107531, 
    0.001107531, 0.001107529, 0.001107529, 0.001107529, 0.001107528, 
    0.001107528, 0.001107526, 0.001107525, 0.001107524, 0.001107524, 
    0.001107524, 0.001107524, 0.001107525, 0.001107524, 0.001107524, 
    0.001107524, 0.001107523, 0.001107523, 0.001107523, 0.001107523, 
    0.00110753, 0.00110753, 0.00110753, 0.00110753, 0.00110753, 0.001107529, 
    0.001107529, 0.001107527, 0.001107528, 0.001107526, 0.001107527, 
    0.001107527, 0.001107526, 0.001107527, 0.001107525, 0.001107527, 
    0.001107524, 0.001107526, 0.001107524, 0.001107524, 0.001107524, 
    0.001107523, 0.001107523, 0.001107522, 0.001107522, 0.001107521, 
    0.001107529, 0.001107529, 0.001107529, 0.001107528, 0.001107528, 
    0.001107527, 0.001107526, 0.001107526, 0.001107526, 0.001107525, 
    0.001107527, 0.001107526, 0.001107529, 0.001107528, 0.001107528, 
    0.001107529, 0.001107526, 0.001107528, 0.001107525, 0.001107526, 
    0.001107523, 0.001107525, 0.001107522, 0.001107521, 0.00110752, 
    0.001107519, 0.001107529, 0.001107529, 0.001107528, 0.001107528, 
    0.001107527, 0.001107526, 0.001107526, 0.001107526, 0.001107525, 
    0.001107525, 0.001107526, 0.001107525, 0.001107528, 0.001107526, 
    0.001107529, 0.001107528, 0.001107528, 0.001107528, 0.001107527, 
    0.001107526, 0.001107525, 0.001107526, 0.001107522, 0.001107523, 
    0.001107518, 0.00110752, 0.001107529, 0.001107529, 0.001107527, 
    0.001107528, 0.001107526, 0.001107525, 0.001107525, 0.001107524, 
    0.001107524, 0.001107524, 0.001107524, 0.001107524, 0.001107526, 
    0.001107525, 0.001107527, 0.001107527, 0.001107527, 0.001107527, 
    0.001107526, 0.001107526, 0.001107525, 0.001107525, 0.001107524, 
    0.001107526, 0.001107521, 0.001107524, 0.001107528, 0.001107527, 
    0.001107527, 0.001107528, 0.001107525, 0.001107526, 0.001107524, 
    0.001107524, 0.001107524, 0.001107524, 0.001107524, 0.001107525, 
    0.001107525, 0.001107526, 0.001107527, 0.001107528, 0.001107527, 
    0.001107527, 0.001107525, 0.001107524, 0.001107524, 0.001107524, 
    0.001107526, 0.001107525, 0.001107525, 0.001107524, 0.001107526, 
    0.001107525, 0.001107527, 0.001107527, 0.001107526, 0.001107525, 
    0.001107525, 0.001107524, 0.001107524, 0.001107525, 0.001107526, 
    0.001107526, 0.001107526, 0.001107527, 0.001107527, 0.001107527, 
    0.001107526, 0.001107525, 0.001107524, 0.001107523, 0.001107523, 
    0.001107522, 0.001107523, 0.001107521, 0.001107523, 0.00110752, 
    0.001107525, 0.001107523, 0.001107526, 0.001107526, 0.001107525, 
    0.001107524, 0.001107524, 0.001107523, 0.001107526, 0.001107527, 
    0.001107527, 0.001107528, 0.001107527, 0.001107527, 0.001107526, 
    0.001107527, 0.001107525, 0.001107526, 0.001107524, 0.001107523, 
    0.001107521, 0.00110752, 0.001107519, 0.001107519, 0.001107518, 
    0.001107518,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N =
  2.684263e-07, 2.684261e-07, 2.684261e-07, 2.684259e-07, 2.68426e-07, 
    2.684259e-07, 2.684263e-07, 2.684261e-07, 2.684262e-07, 2.684263e-07, 
    2.684255e-07, 2.684259e-07, 2.684251e-07, 2.684253e-07, 2.684247e-07, 
    2.684251e-07, 2.684246e-07, 2.684247e-07, 2.684244e-07, 2.684245e-07, 
    2.684241e-07, 2.684243e-07, 2.684239e-07, 2.684241e-07, 2.684241e-07, 
    2.684243e-07, 2.684258e-07, 2.684255e-07, 2.684258e-07, 2.684258e-07, 
    2.684258e-07, 2.68426e-07, 2.684261e-07, 2.684264e-07, 2.684263e-07, 
    2.684262e-07, 2.684258e-07, 2.684259e-07, 2.684256e-07, 2.684256e-07, 
    2.684252e-07, 2.684254e-07, 2.684248e-07, 2.684249e-07, 2.684245e-07, 
    2.684246e-07, 2.684245e-07, 2.684245e-07, 2.684245e-07, 2.684247e-07, 
    2.684246e-07, 2.684247e-07, 2.684254e-07, 2.684252e-07, 2.684257e-07, 
    2.68426e-07, 2.684263e-07, 2.684264e-07, 2.684264e-07, 2.684264e-07, 
    2.684262e-07, 2.68426e-07, 2.684258e-07, 2.684257e-07, 2.684256e-07, 
    2.684253e-07, 2.684251e-07, 2.684247e-07, 2.684248e-07, 2.684247e-07, 
    2.684246e-07, 2.684244e-07, 2.684245e-07, 2.684244e-07, 2.684247e-07, 
    2.684245e-07, 2.684249e-07, 2.684247e-07, 2.684256e-07, 2.684259e-07, 
    2.68426e-07, 2.684261e-07, 2.684264e-07, 2.684262e-07, 2.684263e-07, 
    2.684261e-07, 2.68426e-07, 2.68426e-07, 2.684257e-07, 2.684258e-07, 
    2.684251e-07, 2.684254e-07, 2.684246e-07, 2.684248e-07, 2.684246e-07, 
    2.684247e-07, 2.684245e-07, 2.684247e-07, 2.684243e-07, 2.684243e-07, 
    2.684243e-07, 2.684241e-07, 2.684247e-07, 2.684245e-07, 2.68426e-07, 
    2.68426e-07, 2.68426e-07, 2.684262e-07, 2.684262e-07, 2.684264e-07, 
    2.684262e-07, 2.684261e-07, 2.68426e-07, 2.684259e-07, 2.684258e-07, 
    2.684256e-07, 2.684253e-07, 2.68425e-07, 2.684248e-07, 2.684246e-07, 
    2.684247e-07, 2.684247e-07, 2.684247e-07, 2.684248e-07, 2.684243e-07, 
    2.684246e-07, 2.684241e-07, 2.684242e-07, 2.684244e-07, 2.684242e-07, 
    2.68426e-07, 2.684261e-07, 2.684263e-07, 2.684261e-07, 2.684264e-07, 
    2.684262e-07, 2.684262e-07, 2.684258e-07, 2.684257e-07, 2.684257e-07, 
    2.684255e-07, 2.684254e-07, 2.684251e-07, 2.684248e-07, 2.684246e-07, 
    2.684246e-07, 2.684246e-07, 2.684245e-07, 2.684247e-07, 2.684245e-07, 
    2.684245e-07, 2.684246e-07, 2.684242e-07, 2.684243e-07, 2.684242e-07, 
    2.684243e-07, 2.68426e-07, 2.68426e-07, 2.68426e-07, 2.684259e-07, 
    2.68426e-07, 2.684257e-07, 2.684256e-07, 2.684252e-07, 2.684254e-07, 
    2.684251e-07, 2.684254e-07, 2.684253e-07, 2.684251e-07, 2.684253e-07, 
    2.684248e-07, 2.684252e-07, 2.684245e-07, 2.684249e-07, 2.684245e-07, 
    2.684246e-07, 2.684245e-07, 2.684244e-07, 2.684243e-07, 2.68424e-07, 
    2.684241e-07, 2.684239e-07, 2.684259e-07, 2.684257e-07, 2.684257e-07, 
    2.684256e-07, 2.684255e-07, 2.684253e-07, 2.68425e-07, 2.684251e-07, 
    2.684249e-07, 2.684249e-07, 2.684252e-07, 2.68425e-07, 2.684257e-07, 
    2.684255e-07, 2.684256e-07, 2.684258e-07, 2.684251e-07, 2.684255e-07, 
    2.684248e-07, 2.68425e-07, 2.684244e-07, 2.684247e-07, 2.684241e-07, 
    2.684239e-07, 2.684236e-07, 2.684234e-07, 2.684257e-07, 2.684257e-07, 
    2.684256e-07, 2.684254e-07, 2.684252e-07, 2.68425e-07, 2.684249e-07, 
    2.684249e-07, 2.684248e-07, 2.684247e-07, 2.684249e-07, 2.684247e-07, 
    2.684255e-07, 2.684251e-07, 2.684258e-07, 2.684256e-07, 2.684254e-07, 
    2.684255e-07, 2.684251e-07, 2.684251e-07, 2.684247e-07, 2.684249e-07, 
    2.684239e-07, 2.684244e-07, 2.684232e-07, 2.684235e-07, 2.684258e-07, 
    2.684257e-07, 2.684253e-07, 2.684255e-07, 2.68425e-07, 2.684248e-07, 
    2.684247e-07, 2.684246e-07, 2.684246e-07, 2.684245e-07, 2.684246e-07, 
    2.684245e-07, 2.68425e-07, 2.684248e-07, 2.684253e-07, 2.684252e-07, 
    2.684253e-07, 2.684253e-07, 2.684251e-07, 2.684249e-07, 2.684249e-07, 
    2.684248e-07, 2.684246e-07, 2.68425e-07, 2.684239e-07, 2.684245e-07, 
    2.684255e-07, 2.684253e-07, 2.684253e-07, 2.684254e-07, 2.684249e-07, 
    2.684251e-07, 2.684245e-07, 2.684247e-07, 2.684244e-07, 2.684245e-07, 
    2.684246e-07, 2.684247e-07, 2.684248e-07, 2.68425e-07, 2.684252e-07, 
    2.684254e-07, 2.684253e-07, 2.684252e-07, 2.684249e-07, 2.684246e-07, 
    2.684247e-07, 2.684244e-07, 2.68425e-07, 2.684248e-07, 2.684249e-07, 
    2.684246e-07, 2.684251e-07, 2.684247e-07, 2.684253e-07, 2.684252e-07, 
    2.684251e-07, 2.684247e-07, 2.684247e-07, 2.684246e-07, 2.684247e-07, 
    2.684249e-07, 2.684249e-07, 2.684251e-07, 2.684251e-07, 2.684252e-07, 
    2.684253e-07, 2.684252e-07, 2.684251e-07, 2.684249e-07, 2.684246e-07, 
    2.684244e-07, 2.684243e-07, 2.68424e-07, 2.684243e-07, 2.684239e-07, 
    2.684242e-07, 2.684236e-07, 2.684247e-07, 2.684242e-07, 2.68425e-07, 
    2.684249e-07, 2.684248e-07, 2.684244e-07, 2.684246e-07, 2.684244e-07, 
    2.684249e-07, 2.684252e-07, 2.684252e-07, 2.684254e-07, 2.684252e-07, 
    2.684253e-07, 2.684251e-07, 2.684252e-07, 2.684249e-07, 2.68425e-07, 
    2.684246e-07, 2.684244e-07, 2.684239e-07, 2.684236e-07, 2.684233e-07, 
    2.684232e-07, 2.684232e-07, 2.684232e-07 ;

 LITR2N_TNDNCY_VERT_TRANS =
  -8.82326e-26, 7.352717e-26, -1.323489e-25, -4.41163e-26, 1.02938e-25, 
    -1.078398e-25, 8.333079e-26, -7.352717e-26, -5.391992e-26, 2.695996e-26, 
    1.225453e-26, -1.715634e-25, -1.470543e-26, 1.691125e-25, 9.803622e-26, 
    -8.82326e-26, 3.431268e-26, -1.372507e-25, 1.323489e-25, 1.56858e-25, 
    -2.941087e-26, -2.205815e-26, 1.911706e-25, -2.450905e-26, -8.578169e-26, 
    -9.803622e-26, 5.637083e-26, 1.740143e-25, 5.637083e-26, 2.941087e-26, 
    -6.372354e-26, 5.391992e-26, 3.921449e-26, 7.842898e-26, -1.200944e-25, 
    1.176435e-25, 3.431268e-26, 1.887197e-25, -6.862535e-26, 4.41163e-26, 
    7.352717e-27, -7.597807e-26, -1.29898e-25, 4.65672e-26, -1.54407e-25, 
    6.372354e-26, 1.151926e-25, 1.593089e-25, -3.431268e-26, -3.186177e-26, 
    -1.911706e-25, -8.087988e-26, -1.617598e-25, 7.352717e-26, -5.391992e-26, 
    -1.495052e-25, -9.068351e-26, 2.695996e-26, 2.058761e-25, -2.32836e-25, 
    -8.333079e-26, -7.352717e-26, 4.41163e-26, 1.519561e-25, 6.127264e-26, 
    8.087988e-26, -6.617445e-26, 7.352717e-27, 1.530638e-41, -4.166539e-26, 
    2.769523e-25, -1.593089e-25, 1.02938e-25, -1.715634e-26, 5.391992e-26, 
    -5.882173e-26, 1.740143e-25, -3.431268e-26, -7.842898e-26, -2.450906e-27, 
    -1.323489e-25, -1.960724e-26, 2.426396e-25, -2.450905e-26, 1.740143e-25, 
    2.450906e-25, -1.470543e-26, -9.803622e-27, -1.274471e-25, 1.200944e-25, 
    -5.637083e-26, 1.887197e-25, 1.004871e-25, 3.676358e-26, 2.254833e-25, 
    -5.882173e-26, 1.127417e-25, -2.695996e-26, -8.82326e-26, 1.740143e-25, 
    -8.578169e-26, -2.303851e-25, 5.882173e-26, -1.691125e-25, 6.372354e-26, 
    -3.284213e-25, 3.921449e-26, -1.151926e-25, 1.530638e-41, -1.666616e-25, 
    1.470543e-26, 8.578169e-26, -2.695996e-26, 6.127264e-26, -8.82326e-26, 
    -1.617598e-25, -1.936215e-25, 5.637083e-26, 2.475414e-25, 1.397016e-25, 
    5.882173e-26, 2.401887e-25, 1.151926e-25, -1.200944e-25, -9.313441e-26, 
    5.882173e-26, 1.421525e-25, -4.41163e-26, 1.127417e-25, -1.372507e-25, 
    -1.838179e-25, -1.02938e-25, 1.715634e-26, 2.622469e-25, -1.936215e-25, 
    1.446034e-25, -4.901811e-27, -4.901811e-27, -1.29898e-25, 4.166539e-26, 
    2.401887e-25, 1.225453e-25, -1.225453e-26, -4.166539e-26, -4.41163e-26, 
    -1.54407e-25, 9.558531e-26, 1.446034e-25, 1.078398e-25, 7.107626e-26, 
    1.004871e-25, 1.078398e-25, -1.715634e-26, 1.127417e-25, 8.087988e-26, 
    1.02938e-25, 1.764652e-25, 2.08327e-25, -1.642107e-25, -1.715634e-26, 
    -2.034252e-25, 6.127264e-26, -1.985233e-25, -1.347998e-25, -9.803622e-27, 
    -1.200944e-25, 1.519561e-25, -1.764652e-25, 6.617445e-26, -4.65672e-26, 
    2.32836e-25, 2.671487e-25, 1.372507e-25, 1.715634e-26, 3.676358e-26, 
    5.882173e-26, -1.249962e-25, -1.985233e-25, 1.715634e-26, 7.352717e-27, 
    1.446034e-25, -1.740143e-25, 8.087988e-26, -7.352717e-27, 2.450906e-27, 
    2.450906e-27, -9.803622e-26, -1.225453e-26, -2.941087e-26, -2.279342e-25, 
    1.225453e-26, 1.397016e-25, -1.960724e-26, -2.352869e-25, -8.333079e-26, 
    1.691125e-25, 5.391992e-26, 2.450906e-27, -1.176435e-25, 1.274471e-25, 
    8.578169e-26, 1.323489e-25, 2.401887e-25, -7.107626e-26, 1.495052e-25, 
    3.431268e-26, -9.803622e-27, 7.352717e-26, -2.671487e-25, -8.578169e-26, 
    2.695996e-25, 7.352717e-27, -8.087988e-26, -8.82326e-26, -7.352717e-27, 
    -2.695996e-26, 2.450905e-26, -9.068351e-26, -1.176435e-25, -8.578169e-26, 
    1.372507e-25, 1.200944e-25, 9.313441e-26, -1.274471e-25, 1.446034e-25, 
    -7.107626e-26, -1.323489e-25, 2.132288e-25, 1.225453e-25, 1.960724e-26, 
    -1.715634e-26, -9.803622e-27, -1.593089e-25, -4.215557e-25, 
    -2.450906e-27, -2.009742e-25, 2.450905e-26, -7.842898e-26, -1.81367e-25, 
    -1.397016e-25, 1.053889e-25, 2.450906e-27, 1.470543e-26, 1.470543e-25, 
    1.151926e-25, 5.637083e-26, 2.377378e-25, -8.578169e-26, 8.087988e-26, 
    -2.475414e-25, -3.406759e-25, 1.446034e-25, -8.578169e-26, -1.666616e-25, 
    -2.769523e-25, 1.421525e-25, -1.421525e-25, 4.166539e-26, -3.676358e-26, 
    -4.901811e-26, -3.553813e-25, -2.695996e-25, 2.916578e-25, 1.151926e-25, 
    9.313441e-26, -7.352717e-27, 1.642107e-25, -2.009742e-25, -4.65672e-26, 
    1.470543e-25, -2.990105e-25, -5.637083e-26, -7.352717e-27, -2.695996e-26, 
    6.372354e-26, -2.205815e-25, -1.764652e-25, 1.151926e-25, 1.862688e-25, 
    -1.078398e-25, 8.578169e-26, -1.274471e-25, 9.803622e-27, 2.818541e-25, 
    2.205815e-26, 1.323489e-25, 2.695996e-26, 1.764652e-25, 2.450906e-27, 
    2.548942e-25, 2.573451e-25, 2.08327e-25, -1.249962e-25, -3.210686e-25, 
    1.887197e-25, -7.352717e-27, -6.127264e-26, 1.347998e-25, 1.421525e-25, 
    -2.058761e-25, -7.352717e-27, -2.573451e-25, 1.495052e-25, -2.107779e-25, 
    -2.794032e-25, 5.637083e-26, 4.901811e-26, -1.151926e-25, -7.352717e-26, 
    7.352717e-26, 2.08327e-25, -8.087988e-26, 7.352717e-27, -1.960724e-25, 
    1.225453e-25, -1.225453e-25, 1.078398e-25, -6.127264e-26, 3.921449e-26, 
    -3.431268e-26, 1.960724e-26, 1.02938e-25, -1.960724e-26, -1.274471e-25, 
    1.470543e-25, -6.617445e-26, 1.421525e-25, -1.54407e-25, -7.352717e-26, 
    5.637083e-26, -7.107626e-26, -4.65672e-26, -1.715634e-26, -5.882173e-26, 
    1.02938e-25, -8.087988e-26, 5.882173e-26, -2.524433e-25,
  2.67625e-32, 2.676247e-32, 2.676247e-32, 2.676245e-32, 2.676247e-32, 
    2.676245e-32, 2.676249e-32, 2.676247e-32, 2.676248e-32, 2.676249e-32, 
    2.676241e-32, 2.676245e-32, 2.676237e-32, 2.676239e-32, 2.676233e-32, 
    2.676237e-32, 2.676232e-32, 2.676233e-32, 2.67623e-32, 2.676231e-32, 
    2.676227e-32, 2.676229e-32, 2.676225e-32, 2.676227e-32, 2.676227e-32, 
    2.676229e-32, 2.676244e-32, 2.676242e-32, 2.676244e-32, 2.676244e-32, 
    2.676244e-32, 2.676247e-32, 2.676248e-32, 2.67625e-32, 2.676249e-32, 
    2.676248e-32, 2.676244e-32, 2.676245e-32, 2.676242e-32, 2.676242e-32, 
    2.676238e-32, 2.67624e-32, 2.676234e-32, 2.676236e-32, 2.676231e-32, 
    2.676232e-32, 2.676231e-32, 2.676231e-32, 2.676231e-32, 2.676233e-32, 
    2.676232e-32, 2.676233e-32, 2.67624e-32, 2.676238e-32, 2.676244e-32, 
    2.676247e-32, 2.676249e-32, 2.676251e-32, 2.67625e-32, 2.67625e-32, 
    2.676248e-32, 2.676246e-32, 2.676244e-32, 2.676243e-32, 2.676242e-32, 
    2.676239e-32, 2.676237e-32, 2.676234e-32, 2.676234e-32, 2.676233e-32, 
    2.676232e-32, 2.67623e-32, 2.676231e-32, 2.67623e-32, 2.676233e-32, 
    2.676231e-32, 2.676235e-32, 2.676234e-32, 2.676242e-32, 2.676245e-32, 
    2.676246e-32, 2.676247e-32, 2.67625e-32, 2.676248e-32, 2.676249e-32, 
    2.676247e-32, 2.676246e-32, 2.676247e-32, 2.676243e-32, 2.676244e-32, 
    2.676237e-32, 2.67624e-32, 2.676232e-32, 2.676234e-32, 2.676232e-32, 
    2.676233e-32, 2.676231e-32, 2.676233e-32, 2.676229e-32, 2.676229e-32, 
    2.676229e-32, 2.676227e-32, 2.676233e-32, 2.676231e-32, 2.676247e-32, 
    2.676247e-32, 2.676246e-32, 2.676248e-32, 2.676248e-32, 2.67625e-32, 
    2.676248e-32, 2.676248e-32, 2.676246e-32, 2.676245e-32, 2.676244e-32, 
    2.676242e-32, 2.676239e-32, 2.676236e-32, 2.676234e-32, 2.676232e-32, 
    2.676233e-32, 2.676233e-32, 2.676234e-32, 2.676234e-32, 2.676229e-32, 
    2.676232e-32, 2.676228e-32, 2.676228e-32, 2.67623e-32, 2.676228e-32, 
    2.676247e-32, 2.676247e-32, 2.676249e-32, 2.676247e-32, 2.67625e-32, 
    2.676249e-32, 2.676248e-32, 2.676244e-32, 2.676244e-32, 2.676243e-32, 
    2.676242e-32, 2.67624e-32, 2.676237e-32, 2.676234e-32, 2.676232e-32, 
    2.676232e-32, 2.676232e-32, 2.676232e-32, 2.676233e-32, 2.676232e-32, 
    2.676231e-32, 2.676232e-32, 2.676228e-32, 2.676229e-32, 2.676228e-32, 
    2.676229e-32, 2.676247e-32, 2.676246e-32, 2.676247e-32, 2.676245e-32, 
    2.676246e-32, 2.676243e-32, 2.676242e-32, 2.676238e-32, 2.67624e-32, 
    2.676237e-32, 2.67624e-32, 2.676239e-32, 2.676237e-32, 2.67624e-32, 
    2.676234e-32, 2.676238e-32, 2.676232e-32, 2.676235e-32, 2.676231e-32, 
    2.676232e-32, 2.676231e-32, 2.67623e-32, 2.676229e-32, 2.676227e-32, 
    2.676227e-32, 2.676225e-32, 2.676244e-32, 2.676243e-32, 2.676244e-32, 
    2.676242e-32, 2.676241e-32, 2.676239e-32, 2.676236e-32, 2.676237e-32, 
    2.676235e-32, 2.676235e-32, 2.676238e-32, 2.676236e-32, 2.676243e-32, 
    2.676242e-32, 2.676242e-32, 2.676244e-32, 2.676237e-32, 2.676241e-32, 
    2.676234e-32, 2.676236e-32, 2.67623e-32, 2.676233e-32, 2.676227e-32, 
    2.676225e-32, 2.676222e-32, 2.67622e-32, 2.676243e-32, 2.676244e-32, 
    2.676242e-32, 2.67624e-32, 2.676238e-32, 2.676236e-32, 2.676236e-32, 
    2.676235e-32, 2.676234e-32, 2.676233e-32, 2.676235e-32, 2.676233e-32, 
    2.676241e-32, 2.676237e-32, 2.676244e-32, 2.676242e-32, 2.67624e-32, 
    2.676241e-32, 2.676238e-32, 2.676237e-32, 2.676234e-32, 2.676235e-32, 
    2.676225e-32, 2.67623e-32, 2.676218e-32, 2.676221e-32, 2.676244e-32, 
    2.676243e-32, 2.676239e-32, 2.676241e-32, 2.676236e-32, 2.676234e-32, 
    2.676234e-32, 2.676232e-32, 2.676232e-32, 2.676231e-32, 2.676232e-32, 
    2.676231e-32, 2.676236e-32, 2.676234e-32, 2.676239e-32, 2.676238e-32, 
    2.676239e-32, 2.676239e-32, 2.676237e-32, 2.676235e-32, 2.676235e-32, 
    2.676234e-32, 2.676232e-32, 2.676236e-32, 2.676225e-32, 2.676232e-32, 
    2.676242e-32, 2.676239e-32, 2.676239e-32, 2.67624e-32, 2.676234e-32, 
    2.676237e-32, 2.676231e-32, 2.676233e-32, 2.67623e-32, 2.676232e-32, 
    2.676232e-32, 2.676233e-32, 2.676234e-32, 2.676237e-32, 2.676238e-32, 
    2.67624e-32, 2.676239e-32, 2.676238e-32, 2.676235e-32, 2.676232e-32, 
    2.676233e-32, 2.676231e-32, 2.676236e-32, 2.676234e-32, 2.676235e-32, 
    2.676232e-32, 2.676237e-32, 2.676233e-32, 2.676239e-32, 2.676238e-32, 
    2.676237e-32, 2.676234e-32, 2.676233e-32, 2.676232e-32, 2.676233e-32, 
    2.676235e-32, 2.676235e-32, 2.676237e-32, 2.676237e-32, 2.676238e-32, 
    2.676239e-32, 2.676238e-32, 2.676237e-32, 2.676235e-32, 2.676232e-32, 
    2.67623e-32, 2.676229e-32, 2.676226e-32, 2.676229e-32, 2.676225e-32, 
    2.676228e-32, 2.676222e-32, 2.676233e-32, 2.676228e-32, 2.676237e-32, 
    2.676236e-32, 2.676234e-32, 2.67623e-32, 2.676232e-32, 2.67623e-32, 
    2.676235e-32, 2.676238e-32, 2.676239e-32, 2.67624e-32, 2.676239e-32, 
    2.676239e-32, 2.676237e-32, 2.676238e-32, 2.676235e-32, 2.676236e-32, 
    2.676232e-32, 2.67623e-32, 2.676225e-32, 2.676222e-32, 2.676219e-32, 
    2.676218e-32, 2.676218e-32, 2.676217e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N_TO_SOIL1N =
  2.947935e-15, 2.955894e-15, 2.954348e-15, 2.960762e-15, 2.957206e-15, 
    2.961404e-15, 2.94955e-15, 2.956209e-15, 2.95196e-15, 2.948653e-15, 
    2.973191e-15, 2.961049e-15, 2.985794e-15, 2.978063e-15, 2.99747e-15, 
    2.98459e-15, 3.000065e-15, 2.997101e-15, 3.006024e-15, 3.003469e-15, 
    3.014864e-15, 3.007203e-15, 3.020769e-15, 3.013037e-15, 3.014246e-15, 
    3.00695e-15, 2.963496e-15, 2.97168e-15, 2.963011e-15, 2.964178e-15, 
    2.963655e-15, 2.957279e-15, 2.954062e-15, 2.947328e-15, 2.948551e-15, 
    2.953498e-15, 2.964703e-15, 2.960903e-15, 2.970482e-15, 2.970266e-15, 
    2.980915e-15, 2.976115e-15, 2.993991e-15, 2.988916e-15, 3.003576e-15, 
    2.999891e-15, 3.003402e-15, 3.002338e-15, 3.003416e-15, 2.998011e-15, 
    3.000327e-15, 2.995571e-15, 2.977014e-15, 2.982472e-15, 2.96618e-15, 
    2.956363e-15, 2.949842e-15, 2.94521e-15, 2.945865e-15, 2.947113e-15, 
    2.953527e-15, 2.959555e-15, 2.964144e-15, 2.967213e-15, 2.970235e-15, 
    2.979369e-15, 2.984205e-15, 2.995015e-15, 2.993067e-15, 2.996369e-15, 
    2.999524e-15, 3.004816e-15, 3.003946e-15, 3.006276e-15, 2.996283e-15, 
    3.002925e-15, 2.991959e-15, 2.994958e-15, 2.971048e-15, 2.961929e-15, 
    2.958042e-15, 2.954645e-15, 2.946368e-15, 2.952085e-15, 2.949831e-15, 
    2.955193e-15, 2.958596e-15, 2.956913e-15, 2.967297e-15, 2.963261e-15, 
    2.984491e-15, 2.975354e-15, 2.999156e-15, 2.993467e-15, 3.00052e-15, 
    2.996922e-15, 3.003084e-15, 2.997539e-15, 3.007143e-15, 3.009232e-15, 
    3.007805e-15, 3.01329e-15, 2.997231e-15, 3.003401e-15, 2.956866e-15, 
    2.95714e-15, 2.95842e-15, 2.952794e-15, 2.95245e-15, 2.947294e-15, 
    2.951883e-15, 2.953836e-15, 2.958794e-15, 2.961724e-15, 2.964509e-15, 
    2.970628e-15, 2.977454e-15, 2.986992e-15, 2.993836e-15, 2.998421e-15, 
    2.995611e-15, 2.998092e-15, 2.995318e-15, 2.994018e-15, 3.008449e-15, 
    3.000348e-15, 3.012501e-15, 3.011829e-15, 3.006331e-15, 3.011905e-15, 
    2.957333e-15, 2.955754e-15, 2.950264e-15, 2.95456e-15, 2.946732e-15, 
    2.951114e-15, 2.953632e-15, 2.963344e-15, 2.965478e-15, 2.967454e-15, 
    2.971356e-15, 2.976361e-15, 2.985131e-15, 2.992754e-15, 2.999708e-15, 
    2.999199e-15, 2.999378e-15, 3.00093e-15, 2.997084e-15, 3.001561e-15, 
    3.002311e-15, 3.000348e-15, 3.011739e-15, 3.008487e-15, 3.011815e-15, 
    3.009698e-15, 2.956267e-15, 2.958925e-15, 2.957489e-15, 2.960189e-15, 
    2.958286e-15, 2.966741e-15, 2.969274e-15, 2.981118e-15, 2.976262e-15, 
    2.983992e-15, 2.977048e-15, 2.978278e-15, 2.98424e-15, 2.977424e-15, 
    2.992332e-15, 2.982225e-15, 3.00099e-15, 2.990906e-15, 3.001622e-15, 
    2.999678e-15, 3.002897e-15, 3.005777e-15, 3.009401e-15, 3.01608e-15, 
    3.014534e-15, 3.020118e-15, 2.962887e-15, 2.96633e-15, 2.966029e-15, 
    2.969632e-15, 2.972295e-15, 2.978067e-15, 2.987312e-15, 2.983837e-15, 
    2.990217e-15, 2.991497e-15, 2.981805e-15, 2.987755e-15, 2.968635e-15, 
    2.971726e-15, 2.969887e-15, 2.963157e-15, 2.984636e-15, 2.97362e-15, 
    2.993949e-15, 2.987993e-15, 3.005366e-15, 2.996729e-15, 3.013683e-15, 
    3.020914e-15, 3.027721e-15, 3.035659e-15, 2.968211e-15, 2.965871e-15, 
    2.970061e-15, 2.97585e-15, 2.981222e-15, 2.988356e-15, 2.989086e-15, 
    2.990421e-15, 2.993879e-15, 2.996785e-15, 2.990842e-15, 2.997514e-15, 
    2.972439e-15, 2.985592e-15, 2.964985e-15, 2.971194e-15, 2.97551e-15, 
    2.973619e-15, 2.98344e-15, 2.985753e-15, 2.99514e-15, 2.990291e-15, 
    3.019129e-15, 3.006383e-15, 3.041702e-15, 3.031849e-15, 2.965053e-15, 
    2.968203e-15, 2.979153e-15, 2.973945e-15, 2.988833e-15, 2.99249e-15, 
    2.995465e-15, 2.999263e-15, 2.999675e-15, 3.001924e-15, 2.998237e-15, 
    3.001779e-15, 2.988371e-15, 2.994365e-15, 2.977904e-15, 2.981913e-15, 
    2.98007e-15, 2.978046e-15, 2.984291e-15, 2.990935e-15, 2.99108e-15, 
    2.993207e-15, 2.999197e-15, 2.988893e-15, 3.020767e-15, 3.001093e-15, 
    2.971636e-15, 2.977693e-15, 2.978561e-15, 2.976215e-15, 2.992125e-15, 
    2.986364e-15, 3.00187e-15, 2.997682e-15, 3.004543e-15, 3.001134e-15, 
    3.000633e-15, 2.996253e-15, 2.993524e-15, 2.986628e-15, 2.981011e-15, 
    2.976556e-15, 2.977592e-15, 2.982486e-15, 2.991342e-15, 2.999711e-15, 
    2.997877e-15, 3.004022e-15, 2.987754e-15, 2.994577e-15, 2.991941e-15, 
    2.998816e-15, 2.983744e-15, 2.996573e-15, 2.98046e-15, 2.981875e-15, 
    2.98625e-15, 2.995038e-15, 2.996986e-15, 2.99906e-15, 2.997781e-15, 
    2.991567e-15, 2.99055e-15, 2.986144e-15, 2.984926e-15, 2.981567e-15, 
    2.978784e-15, 2.981326e-15, 2.983994e-15, 2.991571e-15, 2.998389e-15, 
    3.005818e-15, 3.007636e-15, 3.016297e-15, 3.009243e-15, 3.020876e-15, 
    3.010981e-15, 3.028103e-15, 2.997319e-15, 3.010696e-15, 2.986449e-15, 
    2.989066e-15, 2.993792e-15, 3.00463e-15, 2.998784e-15, 3.005622e-15, 
    2.99051e-15, 2.982653e-15, 2.980622e-15, 2.976826e-15, 2.980709e-15, 
    2.980393e-15, 2.984107e-15, 2.982914e-15, 2.991822e-15, 2.987038e-15, 
    3.000619e-15, 3.005569e-15, 3.019532e-15, 3.028077e-15, 3.036769e-15, 
    3.040601e-15, 3.041767e-15, 3.042255e-15 ;

 LITR2N_vr =
  1.532742e-05, 1.532741e-05, 1.532741e-05, 1.53274e-05, 1.53274e-05, 
    1.53274e-05, 1.532742e-05, 1.53274e-05, 1.532741e-05, 1.532742e-05, 
    1.532737e-05, 1.53274e-05, 1.532735e-05, 1.532736e-05, 1.532732e-05, 
    1.532735e-05, 1.532732e-05, 1.532733e-05, 1.532731e-05, 1.532731e-05, 
    1.532729e-05, 1.532731e-05, 1.532728e-05, 1.53273e-05, 1.532729e-05, 
    1.532731e-05, 1.532739e-05, 1.532738e-05, 1.532739e-05, 1.532739e-05, 
    1.532739e-05, 1.53274e-05, 1.532741e-05, 1.532742e-05, 1.532742e-05, 
    1.532741e-05, 1.532739e-05, 1.53274e-05, 1.532738e-05, 1.532738e-05, 
    1.532736e-05, 1.532737e-05, 1.532733e-05, 1.532734e-05, 1.532731e-05, 
    1.532732e-05, 1.532731e-05, 1.532732e-05, 1.532731e-05, 1.532732e-05, 
    1.532732e-05, 1.532733e-05, 1.532736e-05, 1.532735e-05, 1.532739e-05, 
    1.53274e-05, 1.532742e-05, 1.532743e-05, 1.532742e-05, 1.532742e-05, 
    1.532741e-05, 1.53274e-05, 1.532739e-05, 1.532738e-05, 1.532738e-05, 
    1.532736e-05, 1.532735e-05, 1.532733e-05, 1.532733e-05, 1.532733e-05, 
    1.532732e-05, 1.532731e-05, 1.532731e-05, 1.532731e-05, 1.532733e-05, 
    1.532732e-05, 1.532734e-05, 1.532733e-05, 1.532738e-05, 1.532739e-05, 
    1.53274e-05, 1.532741e-05, 1.532742e-05, 1.532741e-05, 1.532742e-05, 
    1.532741e-05, 1.53274e-05, 1.53274e-05, 1.532738e-05, 1.532739e-05, 
    1.532735e-05, 1.532737e-05, 1.532732e-05, 1.532733e-05, 1.532732e-05, 
    1.532733e-05, 1.532731e-05, 1.532732e-05, 1.532731e-05, 1.53273e-05, 
    1.53273e-05, 1.53273e-05, 1.532733e-05, 1.532731e-05, 1.53274e-05, 
    1.53274e-05, 1.53274e-05, 1.532741e-05, 1.532741e-05, 1.532742e-05, 
    1.532741e-05, 1.532741e-05, 1.53274e-05, 1.53274e-05, 1.532739e-05, 
    1.532738e-05, 1.532736e-05, 1.532735e-05, 1.532733e-05, 1.532732e-05, 
    1.532733e-05, 1.532732e-05, 1.532733e-05, 1.532733e-05, 1.53273e-05, 
    1.532732e-05, 1.53273e-05, 1.53273e-05, 1.532731e-05, 1.53273e-05, 
    1.53274e-05, 1.532741e-05, 1.532742e-05, 1.532741e-05, 1.532742e-05, 
    1.532742e-05, 1.532741e-05, 1.532739e-05, 1.532739e-05, 1.532738e-05, 
    1.532738e-05, 1.532737e-05, 1.532735e-05, 1.532733e-05, 1.532732e-05, 
    1.532732e-05, 1.532732e-05, 1.532732e-05, 1.532733e-05, 1.532732e-05, 
    1.532732e-05, 1.532732e-05, 1.53273e-05, 1.53273e-05, 1.53273e-05, 
    1.53273e-05, 1.53274e-05, 1.53274e-05, 1.53274e-05, 1.53274e-05, 
    1.53274e-05, 1.532738e-05, 1.532738e-05, 1.532736e-05, 1.532737e-05, 
    1.532735e-05, 1.532736e-05, 1.532736e-05, 1.532735e-05, 1.532736e-05, 
    1.532734e-05, 1.532736e-05, 1.532732e-05, 1.532734e-05, 1.532732e-05, 
    1.532732e-05, 1.532732e-05, 1.532731e-05, 1.53273e-05, 1.532729e-05, 
    1.532729e-05, 1.532728e-05, 1.532739e-05, 1.532739e-05, 1.532739e-05, 
    1.532738e-05, 1.532737e-05, 1.532736e-05, 1.532734e-05, 1.532735e-05, 
    1.532734e-05, 1.532734e-05, 1.532736e-05, 1.532734e-05, 1.532738e-05, 
    1.532738e-05, 1.532738e-05, 1.532739e-05, 1.532735e-05, 1.532737e-05, 
    1.532733e-05, 1.532734e-05, 1.532731e-05, 1.532733e-05, 1.532729e-05, 
    1.532728e-05, 1.532727e-05, 1.532725e-05, 1.532738e-05, 1.532739e-05, 
    1.532738e-05, 1.532737e-05, 1.532736e-05, 1.532734e-05, 1.532734e-05, 
    1.532734e-05, 1.532733e-05, 1.532733e-05, 1.532734e-05, 1.532732e-05, 
    1.532737e-05, 1.532735e-05, 1.532739e-05, 1.532738e-05, 1.532737e-05, 
    1.532737e-05, 1.532735e-05, 1.532735e-05, 1.532733e-05, 1.532734e-05, 
    1.532728e-05, 1.532731e-05, 1.532724e-05, 1.532726e-05, 1.532739e-05, 
    1.532738e-05, 1.532736e-05, 1.532737e-05, 1.532734e-05, 1.532734e-05, 
    1.532733e-05, 1.532732e-05, 1.532732e-05, 1.532732e-05, 1.532732e-05, 
    1.532732e-05, 1.532734e-05, 1.532733e-05, 1.532736e-05, 1.532736e-05, 
    1.532736e-05, 1.532736e-05, 1.532735e-05, 1.532734e-05, 1.532734e-05, 
    1.532733e-05, 1.532732e-05, 1.532734e-05, 1.532728e-05, 1.532732e-05, 
    1.532738e-05, 1.532736e-05, 1.532736e-05, 1.532737e-05, 1.532734e-05, 
    1.532735e-05, 1.532732e-05, 1.532732e-05, 1.532731e-05, 1.532732e-05, 
    1.532732e-05, 1.532733e-05, 1.532733e-05, 1.532735e-05, 1.532736e-05, 
    1.532737e-05, 1.532736e-05, 1.532735e-05, 1.532734e-05, 1.532732e-05, 
    1.532732e-05, 1.532731e-05, 1.532734e-05, 1.532733e-05, 1.532734e-05, 
    1.532732e-05, 1.532735e-05, 1.532733e-05, 1.532736e-05, 1.532736e-05, 
    1.532735e-05, 1.532733e-05, 1.532733e-05, 1.532732e-05, 1.532732e-05, 
    1.532734e-05, 1.532734e-05, 1.532735e-05, 1.532735e-05, 1.532736e-05, 
    1.532736e-05, 1.532736e-05, 1.532735e-05, 1.532734e-05, 1.532732e-05, 
    1.532731e-05, 1.532731e-05, 1.532729e-05, 1.53273e-05, 1.532728e-05, 
    1.53273e-05, 1.532727e-05, 1.532733e-05, 1.53273e-05, 1.532735e-05, 
    1.532734e-05, 1.532733e-05, 1.532731e-05, 1.532732e-05, 1.532731e-05, 
    1.532734e-05, 1.532735e-05, 1.532736e-05, 1.532736e-05, 1.532736e-05, 
    1.532736e-05, 1.532735e-05, 1.532735e-05, 1.532734e-05, 1.532735e-05, 
    1.532732e-05, 1.532731e-05, 1.532728e-05, 1.532727e-05, 1.532725e-05, 
    1.532724e-05, 1.532724e-05, 1.532724e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2_HR =
  1.065062e-13, 1.067938e-13, 1.067379e-13, 1.069696e-13, 1.068412e-13, 
    1.069928e-13, 1.065646e-13, 1.068051e-13, 1.066516e-13, 1.065321e-13, 
    1.074187e-13, 1.0698e-13, 1.07874e-13, 1.075947e-13, 1.082958e-13, 
    1.078305e-13, 1.083896e-13, 1.082825e-13, 1.086049e-13, 1.085126e-13, 
    1.089243e-13, 1.086475e-13, 1.091376e-13, 1.088583e-13, 1.089019e-13, 
    1.086383e-13, 1.070684e-13, 1.073641e-13, 1.070509e-13, 1.070931e-13, 
    1.070741e-13, 1.068438e-13, 1.067275e-13, 1.064843e-13, 1.065285e-13, 
    1.067072e-13, 1.07112e-13, 1.069747e-13, 1.073208e-13, 1.07313e-13, 
    1.076977e-13, 1.075243e-13, 1.081701e-13, 1.079868e-13, 1.085164e-13, 
    1.083833e-13, 1.085102e-13, 1.084717e-13, 1.085107e-13, 1.083154e-13, 
    1.083991e-13, 1.082272e-13, 1.075568e-13, 1.07754e-13, 1.071654e-13, 
    1.068107e-13, 1.065751e-13, 1.064077e-13, 1.064314e-13, 1.064765e-13, 
    1.067082e-13, 1.06926e-13, 1.070918e-13, 1.072027e-13, 1.073119e-13, 
    1.076419e-13, 1.078166e-13, 1.082072e-13, 1.081368e-13, 1.082561e-13, 
    1.083701e-13, 1.085613e-13, 1.085298e-13, 1.08614e-13, 1.08253e-13, 
    1.084929e-13, 1.080967e-13, 1.082051e-13, 1.073412e-13, 1.070118e-13, 
    1.068714e-13, 1.067486e-13, 1.064496e-13, 1.066561e-13, 1.065747e-13, 
    1.067684e-13, 1.068914e-13, 1.068306e-13, 1.072057e-13, 1.070599e-13, 
    1.078269e-13, 1.074968e-13, 1.083568e-13, 1.081512e-13, 1.08406e-13, 
    1.082761e-13, 1.084987e-13, 1.082983e-13, 1.086453e-13, 1.087208e-13, 
    1.086692e-13, 1.088674e-13, 1.082872e-13, 1.085101e-13, 1.068289e-13, 
    1.068388e-13, 1.06885e-13, 1.066818e-13, 1.066693e-13, 1.06483e-13, 
    1.066488e-13, 1.067194e-13, 1.068985e-13, 1.070044e-13, 1.07105e-13, 
    1.073261e-13, 1.075727e-13, 1.079173e-13, 1.081646e-13, 1.083302e-13, 
    1.082287e-13, 1.083183e-13, 1.082181e-13, 1.081711e-13, 1.086925e-13, 
    1.083998e-13, 1.088389e-13, 1.088146e-13, 1.08616e-13, 1.088174e-13, 
    1.068457e-13, 1.067887e-13, 1.065903e-13, 1.067456e-13, 1.064627e-13, 
    1.066211e-13, 1.06712e-13, 1.070629e-13, 1.0714e-13, 1.072114e-13, 
    1.073524e-13, 1.075332e-13, 1.078501e-13, 1.081255e-13, 1.083767e-13, 
    1.083583e-13, 1.083648e-13, 1.084209e-13, 1.082819e-13, 1.084437e-13, 
    1.084708e-13, 1.083998e-13, 1.088114e-13, 1.086939e-13, 1.088141e-13, 
    1.087376e-13, 1.068072e-13, 1.069033e-13, 1.068514e-13, 1.069489e-13, 
    1.068802e-13, 1.071856e-13, 1.072772e-13, 1.077051e-13, 1.075296e-13, 
    1.078089e-13, 1.07558e-13, 1.076025e-13, 1.078179e-13, 1.075716e-13, 
    1.081102e-13, 1.077451e-13, 1.08423e-13, 1.080587e-13, 1.084459e-13, 
    1.083756e-13, 1.084919e-13, 1.08596e-13, 1.087269e-13, 1.089682e-13, 
    1.089124e-13, 1.091141e-13, 1.070464e-13, 1.071708e-13, 1.071599e-13, 
    1.072901e-13, 1.073863e-13, 1.075948e-13, 1.079289e-13, 1.078033e-13, 
    1.080338e-13, 1.0808e-13, 1.077299e-13, 1.079449e-13, 1.072541e-13, 
    1.073657e-13, 1.072993e-13, 1.070562e-13, 1.078322e-13, 1.074342e-13, 
    1.081686e-13, 1.079534e-13, 1.085811e-13, 1.082691e-13, 1.088816e-13, 
    1.091429e-13, 1.093888e-13, 1.096756e-13, 1.072387e-13, 1.071542e-13, 
    1.073056e-13, 1.075147e-13, 1.077088e-13, 1.079666e-13, 1.07993e-13, 
    1.080412e-13, 1.081661e-13, 1.082711e-13, 1.080564e-13, 1.082974e-13, 
    1.073915e-13, 1.078667e-13, 1.071222e-13, 1.073465e-13, 1.075024e-13, 
    1.074341e-13, 1.07789e-13, 1.078725e-13, 1.082117e-13, 1.080365e-13, 
    1.090784e-13, 1.086179e-13, 1.098939e-13, 1.095379e-13, 1.071247e-13, 
    1.072385e-13, 1.076341e-13, 1.074459e-13, 1.079838e-13, 1.081159e-13, 
    1.082234e-13, 1.083606e-13, 1.083755e-13, 1.084568e-13, 1.083236e-13, 
    1.084515e-13, 1.079671e-13, 1.081837e-13, 1.07589e-13, 1.077338e-13, 
    1.076672e-13, 1.075941e-13, 1.078197e-13, 1.080597e-13, 1.08065e-13, 
    1.081418e-13, 1.083583e-13, 1.07986e-13, 1.091376e-13, 1.084267e-13, 
    1.073625e-13, 1.075813e-13, 1.076127e-13, 1.075279e-13, 1.081027e-13, 
    1.078946e-13, 1.084548e-13, 1.083035e-13, 1.085514e-13, 1.084282e-13, 
    1.084101e-13, 1.082519e-13, 1.081533e-13, 1.079041e-13, 1.077012e-13, 
    1.075402e-13, 1.075777e-13, 1.077545e-13, 1.080744e-13, 1.083768e-13, 
    1.083106e-13, 1.085326e-13, 1.079448e-13, 1.081913e-13, 1.080961e-13, 
    1.083445e-13, 1.078e-13, 1.082634e-13, 1.076813e-13, 1.077324e-13, 
    1.078905e-13, 1.08208e-13, 1.082784e-13, 1.083533e-13, 1.083071e-13, 
    1.080826e-13, 1.080458e-13, 1.078866e-13, 1.078426e-13, 1.077213e-13, 
    1.076208e-13, 1.077126e-13, 1.07809e-13, 1.080827e-13, 1.08329e-13, 
    1.085975e-13, 1.086631e-13, 1.089761e-13, 1.087212e-13, 1.091415e-13, 
    1.08784e-13, 1.094026e-13, 1.082904e-13, 1.087737e-13, 1.078977e-13, 
    1.079922e-13, 1.08163e-13, 1.085545e-13, 1.083433e-13, 1.085904e-13, 
    1.080444e-13, 1.077605e-13, 1.076872e-13, 1.0755e-13, 1.076903e-13, 
    1.076789e-13, 1.078131e-13, 1.0777e-13, 1.080918e-13, 1.07919e-13, 
    1.084096e-13, 1.085885e-13, 1.090929e-13, 1.094016e-13, 1.097157e-13, 
    1.098541e-13, 1.098963e-13, 1.099139e-13 ;

 LITR3C =
  9.697996e-06, 9.697987e-06, 9.697988e-06, 9.69798e-06, 9.697985e-06, 
    9.697979e-06, 9.697994e-06, 9.697986e-06, 9.697991e-06, 9.697995e-06, 
    9.697965e-06, 9.69798e-06, 9.697949e-06, 9.697959e-06, 9.697936e-06, 
    9.697951e-06, 9.697932e-06, 9.697936e-06, 9.697925e-06, 9.697927e-06, 
    9.697914e-06, 9.697923e-06, 9.697907e-06, 9.697917e-06, 9.697915e-06, 
    9.697924e-06, 9.697977e-06, 9.697967e-06, 9.697977e-06, 9.697976e-06, 
    9.697977e-06, 9.697985e-06, 9.697988e-06, 9.697997e-06, 9.697995e-06, 
    9.697989e-06, 9.697976e-06, 9.69798e-06, 9.697968e-06, 9.697968e-06, 
    9.697956e-06, 9.697961e-06, 9.697939e-06, 9.697946e-06, 9.697927e-06, 
    9.697932e-06, 9.697928e-06, 9.697929e-06, 9.697928e-06, 9.697935e-06, 
    9.697932e-06, 9.697937e-06, 9.69796e-06, 9.697954e-06, 9.697974e-06, 
    9.697986e-06, 9.697994e-06, 9.697999e-06, 9.697998e-06, 9.697997e-06, 
    9.697989e-06, 9.697982e-06, 9.697976e-06, 9.697972e-06, 9.697968e-06, 
    9.697957e-06, 9.697951e-06, 9.697938e-06, 9.69794e-06, 9.697937e-06, 
    9.697933e-06, 9.697927e-06, 9.697927e-06, 9.697925e-06, 9.697937e-06, 
    9.697928e-06, 9.697942e-06, 9.697938e-06, 9.697967e-06, 9.697978e-06, 
    9.697984e-06, 9.697987e-06, 9.697997e-06, 9.697991e-06, 9.697994e-06, 
    9.697987e-06, 9.697983e-06, 9.697985e-06, 9.697972e-06, 9.697977e-06, 
    9.697951e-06, 9.697962e-06, 9.697933e-06, 9.69794e-06, 9.697931e-06, 
    9.697936e-06, 9.697928e-06, 9.697935e-06, 9.697924e-06, 9.697921e-06, 
    9.697923e-06, 9.697916e-06, 9.697936e-06, 9.697928e-06, 9.697985e-06, 
    9.697985e-06, 9.697983e-06, 9.69799e-06, 9.69799e-06, 9.697997e-06, 
    9.697991e-06, 9.697988e-06, 9.697983e-06, 9.697979e-06, 9.697976e-06, 
    9.697968e-06, 9.69796e-06, 9.697948e-06, 9.697939e-06, 9.697934e-06, 
    9.697937e-06, 9.697935e-06, 9.697937e-06, 9.697939e-06, 9.697922e-06, 
    9.697932e-06, 9.697917e-06, 9.697917e-06, 9.697925e-06, 9.697917e-06, 
    9.697985e-06, 9.697987e-06, 9.697993e-06, 9.697987e-06, 9.697997e-06, 
    9.697992e-06, 9.697989e-06, 9.697977e-06, 9.697975e-06, 9.697972e-06, 
    9.697967e-06, 9.697961e-06, 9.69795e-06, 9.697941e-06, 9.697933e-06, 
    9.697933e-06, 9.697933e-06, 9.697931e-06, 9.697936e-06, 9.69793e-06, 
    9.697929e-06, 9.697932e-06, 9.697917e-06, 9.697922e-06, 9.697917e-06, 
    9.69792e-06, 9.697986e-06, 9.697982e-06, 9.697984e-06, 9.697981e-06, 
    9.697983e-06, 9.697973e-06, 9.69797e-06, 9.697956e-06, 9.697961e-06, 
    9.697952e-06, 9.69796e-06, 9.697958e-06, 9.697951e-06, 9.69796e-06, 
    9.697941e-06, 9.697954e-06, 9.697931e-06, 9.697943e-06, 9.69793e-06, 
    9.697933e-06, 9.697928e-06, 9.697925e-06, 9.69792e-06, 9.697913e-06, 
    9.697915e-06, 9.697907e-06, 9.697977e-06, 9.697973e-06, 9.697974e-06, 
    9.697969e-06, 9.697966e-06, 9.697959e-06, 9.697947e-06, 9.697952e-06, 
    9.697944e-06, 9.697943e-06, 9.697955e-06, 9.697947e-06, 9.69797e-06, 
    9.697967e-06, 9.697969e-06, 9.697977e-06, 9.697951e-06, 9.697965e-06, 
    9.697939e-06, 9.697947e-06, 9.697926e-06, 9.697937e-06, 9.697916e-06, 
    9.697907e-06, 9.697898e-06, 9.697888e-06, 9.697971e-06, 9.697974e-06, 
    9.697968e-06, 9.697962e-06, 9.697955e-06, 9.697947e-06, 9.697946e-06, 
    9.697944e-06, 9.697939e-06, 9.697936e-06, 9.697943e-06, 9.697936e-06, 
    9.697966e-06, 9.69795e-06, 9.697975e-06, 9.697967e-06, 9.697962e-06, 
    9.697965e-06, 9.697952e-06, 9.697949e-06, 9.697938e-06, 9.697944e-06, 
    9.697908e-06, 9.697925e-06, 9.697881e-06, 9.697893e-06, 9.697975e-06, 
    9.697971e-06, 9.697957e-06, 9.697964e-06, 9.697946e-06, 9.697941e-06, 
    9.697937e-06, 9.697933e-06, 9.697933e-06, 9.69793e-06, 9.697935e-06, 
    9.69793e-06, 9.697947e-06, 9.697939e-06, 9.697959e-06, 9.697955e-06, 
    9.697957e-06, 9.697959e-06, 9.697951e-06, 9.697943e-06, 9.697943e-06, 
    9.69794e-06, 9.697933e-06, 9.697946e-06, 9.697907e-06, 9.697931e-06, 
    9.697967e-06, 9.697959e-06, 9.697958e-06, 9.697961e-06, 9.697942e-06, 
    9.697949e-06, 9.69793e-06, 9.697935e-06, 9.697927e-06, 9.697931e-06, 
    9.697931e-06, 9.697937e-06, 9.69794e-06, 9.697948e-06, 9.697956e-06, 
    9.697961e-06, 9.697959e-06, 9.697954e-06, 9.697943e-06, 9.697933e-06, 
    9.697935e-06, 9.697927e-06, 9.697947e-06, 9.697938e-06, 9.697942e-06, 
    9.697934e-06, 9.697952e-06, 9.697937e-06, 9.697956e-06, 9.697955e-06, 
    9.697949e-06, 9.697938e-06, 9.697936e-06, 9.697933e-06, 9.697935e-06, 
    9.697943e-06, 9.697944e-06, 9.697949e-06, 9.69795e-06, 9.697955e-06, 
    9.697958e-06, 9.697955e-06, 9.697952e-06, 9.697943e-06, 9.697934e-06, 
    9.697925e-06, 9.697923e-06, 9.697912e-06, 9.697921e-06, 9.697907e-06, 
    9.697918e-06, 9.697897e-06, 9.697936e-06, 9.697919e-06, 9.697948e-06, 
    9.697946e-06, 9.69794e-06, 9.697927e-06, 9.697934e-06, 9.697926e-06, 
    9.697944e-06, 9.697954e-06, 9.697956e-06, 9.69796e-06, 9.697956e-06, 
    9.697957e-06, 9.697952e-06, 9.697953e-06, 9.697942e-06, 9.697948e-06, 
    9.697931e-06, 9.697926e-06, 9.697908e-06, 9.697897e-06, 9.697887e-06, 
    9.697883e-06, 9.697881e-06, 9.69788e-06 ;

 LITR3C_TO_SOIL2C =
  5.325308e-14, 5.339687e-14, 5.336894e-14, 5.34848e-14, 5.342056e-14, 
    5.34964e-14, 5.328226e-14, 5.340256e-14, 5.332579e-14, 5.326606e-14, 
    5.370932e-14, 5.348997e-14, 5.393699e-14, 5.379734e-14, 5.41479e-14, 
    5.391524e-14, 5.419478e-14, 5.414124e-14, 5.430243e-14, 5.425628e-14, 
    5.446213e-14, 5.432373e-14, 5.456879e-14, 5.442912e-14, 5.445096e-14, 
    5.431915e-14, 5.353419e-14, 5.368202e-14, 5.352542e-14, 5.354651e-14, 
    5.353706e-14, 5.342187e-14, 5.336376e-14, 5.324212e-14, 5.326421e-14, 
    5.335357e-14, 5.3556e-14, 5.348735e-14, 5.366039e-14, 5.365648e-14, 
    5.384884e-14, 5.376214e-14, 5.408506e-14, 5.399339e-14, 5.425821e-14, 
    5.419164e-14, 5.425507e-14, 5.423584e-14, 5.425532e-14, 5.415769e-14, 
    5.419952e-14, 5.411359e-14, 5.377838e-14, 5.387698e-14, 5.358267e-14, 
    5.340533e-14, 5.328753e-14, 5.320385e-14, 5.321568e-14, 5.323823e-14, 
    5.335409e-14, 5.346298e-14, 5.35459e-14, 5.360133e-14, 5.365592e-14, 
    5.382092e-14, 5.390828e-14, 5.410357e-14, 5.406838e-14, 5.412801e-14, 
    5.418502e-14, 5.428062e-14, 5.426489e-14, 5.430698e-14, 5.412647e-14, 
    5.424645e-14, 5.404835e-14, 5.410254e-14, 5.36706e-14, 5.350588e-14, 
    5.343567e-14, 5.33743e-14, 5.322478e-14, 5.332804e-14, 5.328734e-14, 
    5.338419e-14, 5.344567e-14, 5.341527e-14, 5.360284e-14, 5.352994e-14, 
    5.391346e-14, 5.37484e-14, 5.417837e-14, 5.407561e-14, 5.4203e-14, 
    5.413802e-14, 5.424933e-14, 5.414915e-14, 5.432266e-14, 5.436039e-14, 
    5.43346e-14, 5.443368e-14, 5.414359e-14, 5.425506e-14, 5.341442e-14, 
    5.341937e-14, 5.344248e-14, 5.334086e-14, 5.333465e-14, 5.32415e-14, 
    5.33244e-14, 5.335968e-14, 5.344925e-14, 5.350217e-14, 5.355248e-14, 
    5.366301e-14, 5.378633e-14, 5.395862e-14, 5.408227e-14, 5.41651e-14, 
    5.411433e-14, 5.415915e-14, 5.410903e-14, 5.408554e-14, 5.434624e-14, 
    5.41999e-14, 5.441944e-14, 5.44073e-14, 5.430797e-14, 5.440867e-14, 
    5.342286e-14, 5.339432e-14, 5.329516e-14, 5.337277e-14, 5.323136e-14, 
    5.331051e-14, 5.335599e-14, 5.353143e-14, 5.356999e-14, 5.360568e-14, 
    5.367618e-14, 5.376658e-14, 5.392502e-14, 5.406271e-14, 5.418834e-14, 
    5.417914e-14, 5.418238e-14, 5.421041e-14, 5.414094e-14, 5.422182e-14, 
    5.423537e-14, 5.419991e-14, 5.440568e-14, 5.434693e-14, 5.440705e-14, 
    5.43688e-14, 5.34036e-14, 5.345161e-14, 5.342567e-14, 5.347445e-14, 
    5.344007e-14, 5.359281e-14, 5.363856e-14, 5.385252e-14, 5.376479e-14, 
    5.390443e-14, 5.3779e-14, 5.380122e-14, 5.390892e-14, 5.378579e-14, 
    5.405509e-14, 5.387252e-14, 5.42115e-14, 5.402933e-14, 5.422291e-14, 
    5.41878e-14, 5.424594e-14, 5.429798e-14, 5.436344e-14, 5.448409e-14, 
    5.445617e-14, 5.455704e-14, 5.352318e-14, 5.358538e-14, 5.357994e-14, 
    5.364503e-14, 5.369314e-14, 5.37974e-14, 5.396441e-14, 5.390164e-14, 
    5.401689e-14, 5.404e-14, 5.386492e-14, 5.397242e-14, 5.362702e-14, 
    5.368285e-14, 5.364964e-14, 5.352807e-14, 5.391607e-14, 5.371706e-14, 
    5.408431e-14, 5.397671e-14, 5.429055e-14, 5.413452e-14, 5.444079e-14, 
    5.457142e-14, 5.469439e-14, 5.483777e-14, 5.361935e-14, 5.357709e-14, 
    5.365277e-14, 5.375736e-14, 5.38544e-14, 5.398327e-14, 5.399646e-14, 
    5.402058e-14, 5.408304e-14, 5.413554e-14, 5.402818e-14, 5.41487e-14, 
    5.369574e-14, 5.393334e-14, 5.356109e-14, 5.367325e-14, 5.375121e-14, 
    5.371704e-14, 5.389447e-14, 5.393625e-14, 5.410582e-14, 5.401822e-14, 
    5.453916e-14, 5.430892e-14, 5.494694e-14, 5.476894e-14, 5.356232e-14, 
    5.361922e-14, 5.381702e-14, 5.372295e-14, 5.399188e-14, 5.405795e-14, 
    5.411169e-14, 5.418031e-14, 5.418774e-14, 5.422837e-14, 5.416177e-14, 
    5.422576e-14, 5.398354e-14, 5.409183e-14, 5.379446e-14, 5.386689e-14, 
    5.383359e-14, 5.379702e-14, 5.390983e-14, 5.402986e-14, 5.403247e-14, 
    5.40709e-14, 5.417911e-14, 5.399297e-14, 5.456876e-14, 5.421336e-14, 
    5.368124e-14, 5.379065e-14, 5.380633e-14, 5.376395e-14, 5.405136e-14, 
    5.394728e-14, 5.422739e-14, 5.415175e-14, 5.427568e-14, 5.42141e-14, 
    5.420504e-14, 5.412592e-14, 5.407663e-14, 5.395205e-14, 5.385059e-14, 
    5.377011e-14, 5.378882e-14, 5.387722e-14, 5.403721e-14, 5.418839e-14, 
    5.415527e-14, 5.426626e-14, 5.39724e-14, 5.409566e-14, 5.404803e-14, 
    5.417223e-14, 5.389996e-14, 5.41317e-14, 5.384064e-14, 5.38662e-14, 
    5.394522e-14, 5.410398e-14, 5.413916e-14, 5.417663e-14, 5.415352e-14, 
    5.404127e-14, 5.402289e-14, 5.394331e-14, 5.39213e-14, 5.386064e-14, 
    5.381036e-14, 5.385628e-14, 5.390448e-14, 5.404135e-14, 5.416451e-14, 
    5.429871e-14, 5.433155e-14, 5.448801e-14, 5.436059e-14, 5.457072e-14, 
    5.439199e-14, 5.470129e-14, 5.414519e-14, 5.438683e-14, 5.394883e-14, 
    5.39961e-14, 5.408147e-14, 5.427726e-14, 5.417165e-14, 5.429517e-14, 
    5.402218e-14, 5.388025e-14, 5.384356e-14, 5.377499e-14, 5.384513e-14, 
    5.383943e-14, 5.390651e-14, 5.388496e-14, 5.404589e-14, 5.395947e-14, 
    5.42048e-14, 5.429421e-14, 5.454645e-14, 5.470081e-14, 5.485782e-14, 
    5.492705e-14, 5.494812e-14, 5.495692e-14 ;

 LITR3C_vr =
  0.0005537656, 0.000553765, 0.0005537652, 0.0005537647, 0.0005537649, 
    0.0005537646, 0.0005537655, 0.000553765, 0.0005537653, 0.0005537656, 
    0.0005537638, 0.0005537647, 0.0005537629, 0.0005537635, 0.0005537621, 
    0.000553763, 0.000553762, 0.0005537621, 0.0005537616, 0.0005537617, 
    0.0005537609, 0.0005537614, 0.0005537605, 0.000553761, 0.000553761, 
    0.0005537614, 0.0005537645, 0.0005537639, 0.0005537645, 0.0005537645, 
    0.0005537645, 0.0005537649, 0.0005537652, 0.0005537656, 0.0005537656, 
    0.0005537652, 0.0005537644, 0.0005537647, 0.000553764, 0.0005537641, 
    0.0005537633, 0.0005537636, 0.0005537624, 0.0005537627, 0.0005537617, 
    0.000553762, 0.0005537617, 0.0005537618, 0.0005537617, 0.0005537621, 
    0.0005537619, 0.0005537622, 0.0005537635, 0.0005537632, 0.0005537643, 
    0.000553765, 0.0005537655, 0.0005537658, 0.0005537657, 0.0005537656, 
    0.0005537652, 0.0005537648, 0.0005537645, 0.0005537642, 0.0005537641, 
    0.0005537634, 0.0005537631, 0.0005537623, 0.0005537624, 0.0005537622, 
    0.000553762, 0.0005537616, 0.0005537617, 0.0005537615, 0.0005537622, 
    0.0005537617, 0.0005537625, 0.0005537623, 0.000553764, 0.0005537646, 
    0.0005537649, 0.0005537651, 0.0005537657, 0.0005537653, 0.0005537655, 
    0.0005537651, 0.0005537649, 0.000553765, 0.0005537642, 0.0005537645, 
    0.000553763, 0.0005537636, 0.000553762, 0.0005537624, 0.0005537619, 
    0.0005537621, 0.0005537617, 0.0005537621, 0.0005537614, 0.0005537613, 
    0.0005537614, 0.000553761, 0.0005537621, 0.0005537617, 0.000553765, 
    0.0005537649, 0.0005537649, 0.0005537653, 0.0005537653, 0.0005537656, 
    0.0005537653, 0.0005537652, 0.0005537648, 0.0005537646, 0.0005537644, 
    0.000553764, 0.0005537635, 0.0005537628, 0.0005537624, 0.0005537621, 
    0.0005537622, 0.0005537621, 0.0005537622, 0.0005537624, 0.0005537614, 
    0.0005537619, 0.0005537611, 0.0005537611, 0.0005537615, 0.0005537611, 
    0.0005537649, 0.000553765, 0.0005537655, 0.0005537651, 0.0005537657, 
    0.0005537654, 0.0005537652, 0.0005537645, 0.0005537643, 0.0005537642, 
    0.0005537639, 0.0005537636, 0.000553763, 0.0005537625, 0.000553762, 
    0.000553762, 0.000553762, 0.0005537619, 0.0005537621, 0.0005537618, 
    0.0005537618, 0.0005537619, 0.0005537611, 0.0005537614, 0.0005537611, 
    0.0005537613, 0.000553765, 0.0005537648, 0.0005537649, 0.0005537648, 
    0.0005537649, 0.0005537643, 0.0005537641, 0.0005537632, 0.0005537636, 
    0.0005537631, 0.0005537635, 0.0005537635, 0.0005537631, 0.0005537635, 
    0.0005537625, 0.0005537632, 0.0005537619, 0.0005537626, 0.0005537618, 
    0.000553762, 0.0005537617, 0.0005537616, 0.0005537613, 0.0005537608, 
    0.0005537609, 0.0005537606, 0.0005537645, 0.0005537643, 0.0005537643, 
    0.0005537641, 0.0005537639, 0.0005537635, 0.0005537628, 0.0005537631, 
    0.0005537627, 0.0005537625, 0.0005537632, 0.0005537628, 0.0005537641, 
    0.0005537639, 0.0005537641, 0.0005537645, 0.000553763, 0.0005537638, 
    0.0005537624, 0.0005537628, 0.0005537616, 0.0005537622, 0.000553761, 
    0.0005537605, 0.00055376, 0.0005537595, 0.0005537642, 0.0005537643, 
    0.0005537641, 0.0005537636, 0.0005537632, 0.0005537628, 0.0005537627, 
    0.0005537626, 0.0005537624, 0.0005537622, 0.0005537626, 0.0005537621, 
    0.0005537639, 0.0005537629, 0.0005537644, 0.0005537639, 0.0005537636, 
    0.0005537638, 0.0005537631, 0.0005537629, 0.0005537623, 0.0005537626, 
    0.0005537606, 0.0005537615, 0.000553759, 0.0005537597, 0.0005537644, 
    0.0005537642, 0.0005537634, 0.0005537638, 0.0005537627, 0.0005537625, 
    0.0005537622, 0.000553762, 0.000553762, 0.0005537618, 0.0005537621, 
    0.0005537618, 0.0005537628, 0.0005537624, 0.0005537635, 0.0005537632, 
    0.0005537634, 0.0005537635, 0.0005537631, 0.0005537626, 0.0005537626, 
    0.0005537624, 0.000553762, 0.0005537627, 0.0005537605, 0.0005537618, 
    0.0005537639, 0.0005537635, 0.0005537635, 0.0005537636, 0.0005537625, 
    0.0005537629, 0.0005537618, 0.0005537621, 0.0005537616, 0.0005537618, 
    0.0005537619, 0.0005537622, 0.0005537624, 0.0005537629, 0.0005537633, 
    0.0005537636, 0.0005537635, 0.0005537632, 0.0005537625, 0.000553762, 
    0.0005537621, 0.0005537617, 0.0005537628, 0.0005537623, 0.0005537625, 
    0.000553762, 0.0005537631, 0.0005537622, 0.0005537633, 0.0005537632, 
    0.0005537629, 0.0005537623, 0.0005537621, 0.000553762, 0.0005537621, 
    0.0005537625, 0.0005537626, 0.0005537629, 0.000553763, 0.0005537632, 
    0.0005537634, 0.0005537632, 0.0005537631, 0.0005537625, 0.0005537621, 
    0.0005537616, 0.0005537614, 0.0005537608, 0.0005537613, 0.0005537605, 
    0.0005537612, 0.00055376, 0.0005537621, 0.0005537612, 0.0005537629, 
    0.0005537627, 0.0005537624, 0.0005537616, 0.000553762, 0.0005537616, 
    0.0005537626, 0.0005537632, 0.0005537633, 0.0005537636, 0.0005537633, 
    0.0005537633, 0.0005537631, 0.0005537631, 0.0005537625, 0.0005537628, 
    0.0005537619, 0.0005537616, 0.0005537606, 0.00055376, 0.0005537594, 
    0.0005537591, 0.000553759, 0.000553759,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N =
  1.342132e-07, 1.34213e-07, 1.342131e-07, 1.34213e-07, 1.34213e-07, 
    1.342129e-07, 1.342131e-07, 1.34213e-07, 1.342131e-07, 1.342132e-07, 
    1.342127e-07, 1.342129e-07, 1.342125e-07, 1.342127e-07, 1.342123e-07, 
    1.342125e-07, 1.342123e-07, 1.342123e-07, 1.342122e-07, 1.342122e-07, 
    1.34212e-07, 1.342122e-07, 1.342119e-07, 1.342121e-07, 1.34212e-07, 
    1.342122e-07, 1.342129e-07, 1.342128e-07, 1.342129e-07, 1.342129e-07, 
    1.342129e-07, 1.34213e-07, 1.342131e-07, 1.342132e-07, 1.342132e-07, 
    1.342131e-07, 1.342129e-07, 1.34213e-07, 1.342128e-07, 1.342128e-07, 
    1.342126e-07, 1.342127e-07, 1.342124e-07, 1.342125e-07, 1.342122e-07, 
    1.342123e-07, 1.342122e-07, 1.342122e-07, 1.342122e-07, 1.342123e-07, 
    1.342123e-07, 1.342124e-07, 1.342127e-07, 1.342126e-07, 1.342129e-07, 
    1.34213e-07, 1.342131e-07, 1.342132e-07, 1.342132e-07, 1.342132e-07, 
    1.342131e-07, 1.34213e-07, 1.342129e-07, 1.342128e-07, 1.342128e-07, 
    1.342126e-07, 1.342126e-07, 1.342124e-07, 1.342124e-07, 1.342123e-07, 
    1.342123e-07, 1.342122e-07, 1.342122e-07, 1.342122e-07, 1.342123e-07, 
    1.342122e-07, 1.342124e-07, 1.342124e-07, 1.342128e-07, 1.342129e-07, 
    1.34213e-07, 1.342131e-07, 1.342132e-07, 1.342131e-07, 1.342131e-07, 
    1.34213e-07, 1.34213e-07, 1.34213e-07, 1.342128e-07, 1.342129e-07, 
    1.342125e-07, 1.342127e-07, 1.342123e-07, 1.342124e-07, 1.342123e-07, 
    1.342123e-07, 1.342122e-07, 1.342123e-07, 1.342122e-07, 1.342121e-07, 
    1.342122e-07, 1.342121e-07, 1.342123e-07, 1.342122e-07, 1.34213e-07, 
    1.34213e-07, 1.34213e-07, 1.342131e-07, 1.342131e-07, 1.342132e-07, 
    1.342131e-07, 1.342131e-07, 1.34213e-07, 1.342129e-07, 1.342129e-07, 
    1.342128e-07, 1.342127e-07, 1.342125e-07, 1.342124e-07, 1.342123e-07, 
    1.342124e-07, 1.342123e-07, 1.342124e-07, 1.342124e-07, 1.342121e-07, 
    1.342123e-07, 1.342121e-07, 1.342121e-07, 1.342122e-07, 1.342121e-07, 
    1.34213e-07, 1.34213e-07, 1.342131e-07, 1.342131e-07, 1.342132e-07, 
    1.342131e-07, 1.342131e-07, 1.342129e-07, 1.342129e-07, 1.342128e-07, 
    1.342128e-07, 1.342127e-07, 1.342125e-07, 1.342124e-07, 1.342123e-07, 
    1.342123e-07, 1.342123e-07, 1.342123e-07, 1.342123e-07, 1.342123e-07, 
    1.342122e-07, 1.342123e-07, 1.342121e-07, 1.342121e-07, 1.342121e-07, 
    1.342121e-07, 1.34213e-07, 1.34213e-07, 1.34213e-07, 1.34213e-07, 
    1.34213e-07, 1.342129e-07, 1.342128e-07, 1.342126e-07, 1.342127e-07, 
    1.342126e-07, 1.342127e-07, 1.342127e-07, 1.342126e-07, 1.342127e-07, 
    1.342124e-07, 1.342126e-07, 1.342123e-07, 1.342124e-07, 1.342123e-07, 
    1.342123e-07, 1.342122e-07, 1.342122e-07, 1.342121e-07, 1.34212e-07, 
    1.34212e-07, 1.342119e-07, 1.342129e-07, 1.342129e-07, 1.342129e-07, 
    1.342128e-07, 1.342128e-07, 1.342127e-07, 1.342125e-07, 1.342126e-07, 
    1.342125e-07, 1.342124e-07, 1.342126e-07, 1.342125e-07, 1.342128e-07, 
    1.342128e-07, 1.342128e-07, 1.342129e-07, 1.342125e-07, 1.342127e-07, 
    1.342124e-07, 1.342125e-07, 1.342122e-07, 1.342123e-07, 1.342121e-07, 
    1.342119e-07, 1.342118e-07, 1.342117e-07, 1.342128e-07, 1.342129e-07, 
    1.342128e-07, 1.342127e-07, 1.342126e-07, 1.342125e-07, 1.342125e-07, 
    1.342124e-07, 1.342124e-07, 1.342123e-07, 1.342124e-07, 1.342123e-07, 
    1.342128e-07, 1.342125e-07, 1.342129e-07, 1.342128e-07, 1.342127e-07, 
    1.342127e-07, 1.342126e-07, 1.342125e-07, 1.342124e-07, 1.342124e-07, 
    1.34212e-07, 1.342122e-07, 1.342116e-07, 1.342117e-07, 1.342129e-07, 
    1.342128e-07, 1.342126e-07, 1.342127e-07, 1.342125e-07, 1.342124e-07, 
    1.342124e-07, 1.342123e-07, 1.342123e-07, 1.342123e-07, 1.342123e-07, 
    1.342123e-07, 1.342125e-07, 1.342124e-07, 1.342127e-07, 1.342126e-07, 
    1.342126e-07, 1.342127e-07, 1.342126e-07, 1.342124e-07, 1.342124e-07, 
    1.342124e-07, 1.342123e-07, 1.342125e-07, 1.342119e-07, 1.342123e-07, 
    1.342128e-07, 1.342127e-07, 1.342126e-07, 1.342127e-07, 1.342124e-07, 
    1.342125e-07, 1.342123e-07, 1.342123e-07, 1.342122e-07, 1.342123e-07, 
    1.342123e-07, 1.342123e-07, 1.342124e-07, 1.342125e-07, 1.342126e-07, 
    1.342127e-07, 1.342127e-07, 1.342126e-07, 1.342124e-07, 1.342123e-07, 
    1.342123e-07, 1.342122e-07, 1.342125e-07, 1.342124e-07, 1.342124e-07, 
    1.342123e-07, 1.342126e-07, 1.342123e-07, 1.342126e-07, 1.342126e-07, 
    1.342125e-07, 1.342124e-07, 1.342123e-07, 1.342123e-07, 1.342123e-07, 
    1.342124e-07, 1.342124e-07, 1.342125e-07, 1.342125e-07, 1.342126e-07, 
    1.342126e-07, 1.342126e-07, 1.342126e-07, 1.342124e-07, 1.342123e-07, 
    1.342122e-07, 1.342122e-07, 1.34212e-07, 1.342121e-07, 1.342119e-07, 
    1.342121e-07, 1.342118e-07, 1.342123e-07, 1.342121e-07, 1.342125e-07, 
    1.342125e-07, 1.342124e-07, 1.342122e-07, 1.342123e-07, 1.342122e-07, 
    1.342124e-07, 1.342126e-07, 1.342126e-07, 1.342127e-07, 1.342126e-07, 
    1.342126e-07, 1.342126e-07, 1.342126e-07, 1.342124e-07, 1.342125e-07, 
    1.342123e-07, 1.342122e-07, 1.34212e-07, 1.342118e-07, 1.342117e-07, 
    1.342116e-07, 1.342116e-07, 1.342116e-07 ;

 LITR3N_TNDNCY_VERT_TRANS =
  -6.617445e-26, -7.352717e-27, -4.901811e-27, 1.629852e-25, -5.269447e-26, 
    1.078398e-25, 4.534175e-26, -1.225453e-27, 1.225453e-27, -2.941087e-26, 
    -5.024356e-26, -3.676358e-27, -5.391992e-26, -6.98508e-26, -1.004871e-25, 
    3.063632e-26, -1.960724e-26, -4.166539e-26, -1.470543e-26, -1.004871e-25, 
    6.127264e-26, -2.450906e-27, 5.759628e-26, 2.695996e-26, 7.352717e-27, 
    -4.043994e-26, 1.593089e-26, -6.127264e-27, 9.558531e-26, -1.225453e-26, 
    -7.720352e-26, -7.597807e-26, 3.676358e-27, -6.127264e-27, -8.333079e-26, 
    -1.838179e-26, -1.593089e-26, 3.431268e-26, -6.617445e-26, -9.803622e-27, 
    5.759628e-26, 8.578169e-26, 1.838179e-26, -5.882173e-26, -4.289085e-26, 
    6.4949e-26, -5.637083e-26, 8.333079e-26, 4.166539e-26, -3.798904e-26, 
    -5.391992e-26, -6.372354e-26, 6.4949e-26, -7.352717e-27, 1.838179e-26, 
    3.676358e-26, 6.004719e-26, 3.308722e-26, -2.450905e-26, 7.107626e-26, 
    -1.286725e-25, -2.941087e-26, -2.450905e-26, -8.945805e-26, 
    -2.818541e-26, 2.08327e-26, 8.455624e-26, 3.431268e-26, -6.862535e-26, 
    -7.352717e-27, -2.818541e-26, -1.838179e-26, 7.352717e-27, 7.475262e-26, 
    1.102908e-26, 6.249809e-26, 6.127264e-27, -3.921449e-26, -3.063632e-26, 
    2.08327e-26, 1.225453e-26, -7.230172e-26, -6.372354e-26, -1.29898e-25, 
    1.470543e-25, -1.703379e-25, -3.921449e-26, -8.333079e-26, -6.862535e-26, 
    7.107626e-26, -1.102908e-25, 3.676358e-27, -5.637083e-26, 4.901811e-27, 
    4.901811e-27, -2.32836e-26, 2.450906e-27, 1.225453e-26, 1.286725e-25, 
    -9.803622e-27, 1.017126e-25, -7.352717e-27, -5.024356e-26, 4.901811e-26, 
    -4.901811e-27, 4.534175e-26, 1.838179e-26, 3.676358e-26, 6.372354e-26, 
    -6.249809e-26, -9.681077e-26, 3.308722e-26, 8.700715e-26, -4.779266e-26, 
    4.901811e-26, 6.862535e-26, -8.82326e-26, 5.759628e-26, 3.676358e-27, 
    -1.225453e-27, 2.08327e-26, 3.921449e-26, 2.08327e-26, 1.838179e-26, 
    -8.087988e-26, 1.004871e-25, -3.553813e-26, -5.146902e-26, -1.470543e-25, 
    -1.078398e-25, 1.960724e-26, -5.146902e-26, 1.593089e-26, 9.558531e-26, 
    -1.225453e-25, 8.210533e-26, 1.936215e-25, 3.431268e-26, -1.715634e-26, 
    1.347998e-26, -2.450905e-26, -3.063632e-26, 1.225453e-27, 1.409271e-25, 
    8.210533e-26, 2.450905e-26, 7.352717e-27, -2.573451e-26, -3.431268e-26, 
    -4.289085e-26, 8.578169e-27, 2.450905e-26, -6.73999e-26, 1.004871e-25, 
    7.652491e-42, -8.578169e-26, -2.205815e-26, 7.352717e-27, -1.960724e-26, 
    -5.146902e-26, 1.127417e-25, 1.102908e-26, 3.308722e-26, 1.090653e-25, 
    -5.637083e-26, 2.450905e-26, -1.960724e-26, -3.798904e-26, -5.391992e-26, 
    1.838179e-25, 3.676358e-26, -4.289085e-26, -1.16418e-25, -4.65672e-26, 
    9.803622e-27, 6.004719e-26, 9.803622e-27, 1.593089e-26, -4.901811e-27, 
    -1.580834e-25, -2.450906e-27, 2.205815e-26, -1.066144e-25, 4.41163e-26, 
    3.553813e-26, 8.700715e-26, -3.186177e-26, -4.534175e-26, 2.08327e-26, 
    -3.308722e-26, -7.352717e-26, 1.066144e-25, -8.333079e-26, 9.558531e-26, 
    -5.637083e-26, -5.269447e-26, -5.637083e-26, -1.225453e-26, 2.695996e-26, 
    6.862535e-26, -9.558531e-26, 6.004719e-26, -5.269447e-26, 2.941087e-26, 
    8.578169e-27, -5.514538e-26, 2.205815e-26, 1.347998e-26, -1.960724e-26, 
    6.127264e-27, -4.779266e-26, -2.32836e-26, 1.470543e-26, -3.553813e-26, 
    -9.803622e-27, -2.205815e-26, 5.146902e-26, -6.127264e-26, -2.450905e-26, 
    1.225453e-27, 2.818541e-26, 1.225453e-25, -2.450905e-26, -2.573451e-26, 
    -4.166539e-26, 2.08327e-26, 8.333079e-26, -1.115162e-25, -2.205815e-26, 
    -1.004871e-25, -1.43378e-25, 0, -3.308722e-26, 7.352717e-27, 
    1.176435e-25, 8.333079e-26, -2.818541e-26, 9.558531e-26, 6.73999e-26, 
    -1.004871e-25, -1.960724e-26, -7.107626e-26, -2.205815e-26, -8.82326e-26, 
    5.146902e-26, 1.102908e-26, -1.225453e-27, 2.573451e-26, 4.41163e-26, 
    -2.450906e-27, -4.043994e-26, 2.32836e-26, 2.941087e-26, -1.225453e-27, 
    7.652491e-42, 2.818541e-26, 1.838179e-26, -1.102908e-26, -6.127264e-27, 
    -7.352717e-27, -1.715634e-26, -5.146902e-26, -1.017126e-25, 6.4949e-26, 
    -1.225453e-27, 5.882173e-26, 3.308722e-26, -3.553813e-26, 4.779266e-26, 
    -2.818541e-26, -8.578169e-27, -7.230172e-26, -7.230172e-26, 1.531816e-25, 
    -3.553813e-26, 6.4949e-26, -9.558531e-26, 5.024356e-26, 6.862535e-26, 
    -2.205815e-26, -1.066144e-25, -1.470543e-26, 3.063632e-26, -5.759628e-26, 
    5.024356e-26, 6.004719e-26, -2.450905e-26, -2.450905e-26, 5.391992e-26, 
    3.676358e-27, -4.166539e-26, 7.965443e-26, -7.352717e-26, -2.941087e-26, 
    -5.146902e-26, 1.102908e-26, -1.593089e-26, 2.205815e-26, 1.470543e-26, 
    -6.617445e-26, 3.186177e-26, 3.676358e-26, 4.41163e-26, 6.372354e-26, 
    -6.372354e-26, 4.41163e-26, 8.333079e-26, 1.347998e-26, -3.063632e-26, 
    -7.475262e-26, -4.41163e-26, -1.262216e-25, 4.901811e-27, -7.352717e-26, 
    2.205815e-26, -4.043994e-26, 3.063632e-26, 5.514538e-26, -1.470543e-25, 
    1.56858e-25, 4.65672e-26, 2.450906e-27, 3.676358e-27, -3.676358e-27, 
    1.066144e-25, -1.838179e-26, 1.017126e-25, 6.4949e-26, -6.98508e-26, 
    2.205815e-26, 5.637083e-26, 1.041635e-25, 3.186177e-26, 2.450906e-27, 
    8.578169e-27, -1.225453e-25, -4.901811e-26, 2.818541e-26,
  1.338125e-32, 1.338123e-32, 1.338124e-32, 1.338123e-32, 1.338123e-32, 
    1.338123e-32, 1.338124e-32, 1.338123e-32, 1.338124e-32, 1.338125e-32, 
    1.33812e-32, 1.338123e-32, 1.338118e-32, 1.33812e-32, 1.338116e-32, 
    1.338119e-32, 1.338116e-32, 1.338116e-32, 1.338115e-32, 1.338115e-32, 
    1.338113e-32, 1.338115e-32, 1.338112e-32, 1.338114e-32, 1.338113e-32, 
    1.338115e-32, 1.338122e-32, 1.338121e-32, 1.338122e-32, 1.338122e-32, 
    1.338122e-32, 1.338123e-32, 1.338124e-32, 1.338125e-32, 1.338125e-32, 
    1.338124e-32, 1.338122e-32, 1.338123e-32, 1.338121e-32, 1.338121e-32, 
    1.338119e-32, 1.33812e-32, 1.338117e-32, 1.338118e-32, 1.338115e-32, 
    1.338116e-32, 1.338115e-32, 1.338115e-32, 1.338115e-32, 1.338116e-32, 
    1.338116e-32, 1.338117e-32, 1.33812e-32, 1.338119e-32, 1.338122e-32, 
    1.338123e-32, 1.338124e-32, 1.338125e-32, 1.338125e-32, 1.338125e-32, 
    1.338124e-32, 1.338123e-32, 1.338122e-32, 1.338121e-32, 1.338121e-32, 
    1.338119e-32, 1.338119e-32, 1.338117e-32, 1.338117e-32, 1.338117e-32, 
    1.338116e-32, 1.338115e-32, 1.338115e-32, 1.338115e-32, 1.338117e-32, 
    1.338115e-32, 1.338117e-32, 1.338117e-32, 1.338121e-32, 1.338122e-32, 
    1.338123e-32, 1.338124e-32, 1.338125e-32, 1.338124e-32, 1.338124e-32, 
    1.338124e-32, 1.338123e-32, 1.338123e-32, 1.338121e-32, 1.338122e-32, 
    1.338119e-32, 1.33812e-32, 1.338116e-32, 1.338117e-32, 1.338116e-32, 
    1.338116e-32, 1.338115e-32, 1.338116e-32, 1.338115e-32, 1.338114e-32, 
    1.338115e-32, 1.338114e-32, 1.338116e-32, 1.338115e-32, 1.338123e-32, 
    1.338123e-32, 1.338123e-32, 1.338124e-32, 1.338124e-32, 1.338125e-32, 
    1.338124e-32, 1.338124e-32, 1.338123e-32, 1.338122e-32, 1.338122e-32, 
    1.338121e-32, 1.33812e-32, 1.338118e-32, 1.338117e-32, 1.338116e-32, 
    1.338117e-32, 1.338116e-32, 1.338117e-32, 1.338117e-32, 1.338114e-32, 
    1.338116e-32, 1.338114e-32, 1.338114e-32, 1.338115e-32, 1.338114e-32, 
    1.338123e-32, 1.338123e-32, 1.338124e-32, 1.338124e-32, 1.338125e-32, 
    1.338124e-32, 1.338124e-32, 1.338122e-32, 1.338122e-32, 1.338121e-32, 
    1.338121e-32, 1.33812e-32, 1.338118e-32, 1.338117e-32, 1.338116e-32, 
    1.338116e-32, 1.338116e-32, 1.338116e-32, 1.338116e-32, 1.338116e-32, 
    1.338115e-32, 1.338116e-32, 1.338114e-32, 1.338114e-32, 1.338114e-32, 
    1.338114e-32, 1.338123e-32, 1.338123e-32, 1.338123e-32, 1.338123e-32, 
    1.338123e-32, 1.338121e-32, 1.338121e-32, 1.338119e-32, 1.33812e-32, 
    1.338119e-32, 1.33812e-32, 1.33812e-32, 1.338119e-32, 1.33812e-32, 
    1.338117e-32, 1.338119e-32, 1.338116e-32, 1.338117e-32, 1.338116e-32, 
    1.338116e-32, 1.338115e-32, 1.338115e-32, 1.338114e-32, 1.338113e-32, 
    1.338113e-32, 1.338113e-32, 1.338122e-32, 1.338122e-32, 1.338122e-32, 
    1.338121e-32, 1.338121e-32, 1.33812e-32, 1.338118e-32, 1.338119e-32, 
    1.338118e-32, 1.338117e-32, 1.338119e-32, 1.338118e-32, 1.338121e-32, 
    1.338121e-32, 1.338121e-32, 1.338122e-32, 1.338119e-32, 1.33812e-32, 
    1.338117e-32, 1.338118e-32, 1.338115e-32, 1.338117e-32, 1.338114e-32, 
    1.338112e-32, 1.338111e-32, 1.33811e-32, 1.338121e-32, 1.338122e-32, 
    1.338121e-32, 1.33812e-32, 1.338119e-32, 1.338118e-32, 1.338118e-32, 
    1.338118e-32, 1.338117e-32, 1.338117e-32, 1.338118e-32, 1.338116e-32, 
    1.338121e-32, 1.338118e-32, 1.338122e-32, 1.338121e-32, 1.33812e-32, 
    1.33812e-32, 1.338119e-32, 1.338118e-32, 1.338117e-32, 1.338118e-32, 
    1.338113e-32, 1.338115e-32, 1.338109e-32, 1.33811e-32, 1.338122e-32, 
    1.338121e-32, 1.338119e-32, 1.33812e-32, 1.338118e-32, 1.338117e-32, 
    1.338117e-32, 1.338116e-32, 1.338116e-32, 1.338116e-32, 1.338116e-32, 
    1.338116e-32, 1.338118e-32, 1.338117e-32, 1.33812e-32, 1.338119e-32, 
    1.338119e-32, 1.33812e-32, 1.338119e-32, 1.338117e-32, 1.338117e-32, 
    1.338117e-32, 1.338116e-32, 1.338118e-32, 1.338112e-32, 1.338116e-32, 
    1.338121e-32, 1.33812e-32, 1.33812e-32, 1.33812e-32, 1.338117e-32, 
    1.338118e-32, 1.338116e-32, 1.338116e-32, 1.338115e-32, 1.338116e-32, 
    1.338116e-32, 1.338117e-32, 1.338117e-32, 1.338118e-32, 1.338119e-32, 
    1.33812e-32, 1.33812e-32, 1.338119e-32, 1.338117e-32, 1.338116e-32, 
    1.338116e-32, 1.338115e-32, 1.338118e-32, 1.338117e-32, 1.338117e-32, 
    1.338116e-32, 1.338119e-32, 1.338117e-32, 1.338119e-32, 1.338119e-32, 
    1.338118e-32, 1.338117e-32, 1.338116e-32, 1.338116e-32, 1.338116e-32, 
    1.338117e-32, 1.338118e-32, 1.338118e-32, 1.338118e-32, 1.338119e-32, 
    1.33812e-32, 1.338119e-32, 1.338119e-32, 1.338117e-32, 1.338116e-32, 
    1.338115e-32, 1.338115e-32, 1.338113e-32, 1.338114e-32, 1.338112e-32, 
    1.338114e-32, 1.338111e-32, 1.338116e-32, 1.338114e-32, 1.338118e-32, 
    1.338118e-32, 1.338117e-32, 1.338115e-32, 1.338116e-32, 1.338115e-32, 
    1.338118e-32, 1.338119e-32, 1.338119e-32, 1.33812e-32, 1.338119e-32, 
    1.338119e-32, 1.338119e-32, 1.338119e-32, 1.338117e-32, 1.338118e-32, 
    1.338116e-32, 1.338115e-32, 1.338113e-32, 1.338111e-32, 1.33811e-32, 
    1.338109e-32, 1.338109e-32, 1.338109e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N_TO_SOIL2N =
  1.473967e-15, 1.477947e-15, 1.477174e-15, 1.480381e-15, 1.478603e-15, 
    1.480702e-15, 1.474775e-15, 1.478105e-15, 1.47598e-15, 1.474327e-15, 
    1.486596e-15, 1.480524e-15, 1.492897e-15, 1.489032e-15, 1.498735e-15, 
    1.492295e-15, 1.500032e-15, 1.49855e-15, 1.503012e-15, 1.501734e-15, 
    1.507432e-15, 1.503601e-15, 1.510384e-15, 1.506518e-15, 1.507123e-15, 
    1.503475e-15, 1.481748e-15, 1.48584e-15, 1.481505e-15, 1.482089e-15, 
    1.481827e-15, 1.478639e-15, 1.477031e-15, 1.473664e-15, 1.474276e-15, 
    1.476749e-15, 1.482352e-15, 1.480451e-15, 1.485241e-15, 1.485133e-15, 
    1.490457e-15, 1.488058e-15, 1.496995e-15, 1.494458e-15, 1.501788e-15, 
    1.499945e-15, 1.501701e-15, 1.501169e-15, 1.501708e-15, 1.499006e-15, 
    1.500164e-15, 1.497785e-15, 1.488507e-15, 1.491236e-15, 1.48309e-15, 
    1.478181e-15, 1.474921e-15, 1.472605e-15, 1.472932e-15, 1.473556e-15, 
    1.476763e-15, 1.479777e-15, 1.482072e-15, 1.483606e-15, 1.485117e-15, 
    1.489684e-15, 1.492102e-15, 1.497508e-15, 1.496534e-15, 1.498184e-15, 
    1.499762e-15, 1.502408e-15, 1.501973e-15, 1.503138e-15, 1.498142e-15, 
    1.501462e-15, 1.495979e-15, 1.497479e-15, 1.485524e-15, 1.480964e-15, 
    1.479021e-15, 1.477323e-15, 1.473184e-15, 1.476042e-15, 1.474916e-15, 
    1.477596e-15, 1.479298e-15, 1.478457e-15, 1.483648e-15, 1.481631e-15, 
    1.492246e-15, 1.487677e-15, 1.499578e-15, 1.496734e-15, 1.50026e-15, 
    1.498461e-15, 1.501542e-15, 1.498769e-15, 1.503572e-15, 1.504616e-15, 
    1.503902e-15, 1.506645e-15, 1.498615e-15, 1.501701e-15, 1.478433e-15, 
    1.47857e-15, 1.47921e-15, 1.476397e-15, 1.476225e-15, 1.473647e-15, 
    1.475941e-15, 1.476918e-15, 1.479397e-15, 1.480862e-15, 1.482254e-15, 
    1.485314e-15, 1.488727e-15, 1.493496e-15, 1.496918e-15, 1.499211e-15, 
    1.497805e-15, 1.499046e-15, 1.497659e-15, 1.497009e-15, 1.504224e-15, 
    1.500174e-15, 1.50625e-15, 1.505915e-15, 1.503165e-15, 1.505952e-15, 
    1.478667e-15, 1.477877e-15, 1.475132e-15, 1.47728e-15, 1.473366e-15, 
    1.475557e-15, 1.476816e-15, 1.481672e-15, 1.482739e-15, 1.483727e-15, 
    1.485678e-15, 1.48818e-15, 1.492566e-15, 1.496377e-15, 1.499854e-15, 
    1.4996e-15, 1.499689e-15, 1.500465e-15, 1.498542e-15, 1.500781e-15, 
    1.501156e-15, 1.500174e-15, 1.50587e-15, 1.504243e-15, 1.505907e-15, 
    1.504849e-15, 1.478134e-15, 1.479463e-15, 1.478744e-15, 1.480094e-15, 
    1.479143e-15, 1.48337e-15, 1.484637e-15, 1.490559e-15, 1.488131e-15, 
    1.491996e-15, 1.488524e-15, 1.489139e-15, 1.49212e-15, 1.488712e-15, 
    1.496166e-15, 1.491113e-15, 1.500495e-15, 1.495453e-15, 1.500811e-15, 
    1.499839e-15, 1.501448e-15, 1.502889e-15, 1.5047e-15, 1.50804e-15, 
    1.507267e-15, 1.510059e-15, 1.481443e-15, 1.483165e-15, 1.483014e-15, 
    1.484816e-15, 1.486148e-15, 1.489033e-15, 1.493656e-15, 1.491919e-15, 
    1.495108e-15, 1.495748e-15, 1.490902e-15, 1.493877e-15, 1.484317e-15, 
    1.485863e-15, 1.484943e-15, 1.481579e-15, 1.492318e-15, 1.48681e-15, 
    1.496974e-15, 1.493996e-15, 1.502683e-15, 1.498364e-15, 1.506841e-15, 
    1.510457e-15, 1.513861e-15, 1.517829e-15, 1.484105e-15, 1.482936e-15, 
    1.48503e-15, 1.487925e-15, 1.490611e-15, 1.494178e-15, 1.494543e-15, 
    1.495211e-15, 1.496939e-15, 1.498392e-15, 1.495421e-15, 1.498757e-15, 
    1.486219e-15, 1.492796e-15, 1.482493e-15, 1.485597e-15, 1.487755e-15, 
    1.486809e-15, 1.49172e-15, 1.492876e-15, 1.49757e-15, 1.495145e-15, 
    1.509564e-15, 1.503191e-15, 1.520851e-15, 1.515924e-15, 1.482527e-15, 
    1.484102e-15, 1.489576e-15, 1.486973e-15, 1.494416e-15, 1.496245e-15, 
    1.497733e-15, 1.499632e-15, 1.499837e-15, 1.500962e-15, 1.499119e-15, 
    1.50089e-15, 1.494185e-15, 1.497183e-15, 1.488952e-15, 1.490957e-15, 
    1.490035e-15, 1.489023e-15, 1.492145e-15, 1.495467e-15, 1.49554e-15, 
    1.496603e-15, 1.499599e-15, 1.494446e-15, 1.510383e-15, 1.500546e-15, 
    1.485818e-15, 1.488847e-15, 1.489281e-15, 1.488108e-15, 1.496063e-15, 
    1.493182e-15, 1.500935e-15, 1.498841e-15, 1.502271e-15, 1.500567e-15, 
    1.500316e-15, 1.498126e-15, 1.496762e-15, 1.493314e-15, 1.490506e-15, 
    1.488278e-15, 1.488796e-15, 1.491243e-15, 1.495671e-15, 1.499855e-15, 
    1.498939e-15, 1.502011e-15, 1.493877e-15, 1.497289e-15, 1.495971e-15, 
    1.499408e-15, 1.491872e-15, 1.498286e-15, 1.49023e-15, 1.490937e-15, 
    1.493125e-15, 1.497519e-15, 1.498493e-15, 1.49953e-15, 1.49889e-15, 
    1.495783e-15, 1.495275e-15, 1.493072e-15, 1.492463e-15, 1.490784e-15, 
    1.489392e-15, 1.490663e-15, 1.491997e-15, 1.495785e-15, 1.499194e-15, 
    1.502909e-15, 1.503818e-15, 1.508149e-15, 1.504622e-15, 1.510438e-15, 
    1.505491e-15, 1.514052e-15, 1.49866e-15, 1.505348e-15, 1.493225e-15, 
    1.494533e-15, 1.496896e-15, 1.502315e-15, 1.499392e-15, 1.502811e-15, 
    1.495255e-15, 1.491326e-15, 1.490311e-15, 1.488413e-15, 1.490354e-15, 
    1.490197e-15, 1.492053e-15, 1.491457e-15, 1.495911e-15, 1.493519e-15, 
    1.50031e-15, 1.502784e-15, 1.509766e-15, 1.514038e-15, 1.518384e-15, 
    1.5203e-15, 1.520884e-15, 1.521127e-15 ;

 LITR3N_vr =
  7.663711e-06, 7.663702e-06, 7.663704e-06, 7.663698e-06, 7.663702e-06, 
    7.663697e-06, 7.663709e-06, 7.663702e-06, 7.663707e-06, 7.66371e-06, 
    7.663686e-06, 7.663698e-06, 7.663673e-06, 7.663682e-06, 7.663662e-06, 
    7.663675e-06, 7.66366e-06, 7.663662e-06, 7.663654e-06, 7.663657e-06, 
    7.663646e-06, 7.663653e-06, 7.66364e-06, 7.663647e-06, 7.663646e-06, 
    7.663653e-06, 7.663695e-06, 7.663688e-06, 7.663696e-06, 7.663695e-06, 
    7.663695e-06, 7.663702e-06, 7.663704e-06, 7.663711e-06, 7.66371e-06, 
    7.663705e-06, 7.663694e-06, 7.663698e-06, 7.663689e-06, 7.663689e-06, 
    7.663679e-06, 7.663683e-06, 7.663666e-06, 7.663671e-06, 7.663657e-06, 
    7.66366e-06, 7.663657e-06, 7.663658e-06, 7.663657e-06, 7.663662e-06, 
    7.66366e-06, 7.663664e-06, 7.663682e-06, 7.663677e-06, 7.663692e-06, 
    7.663702e-06, 7.663709e-06, 7.663713e-06, 7.663712e-06, 7.663712e-06, 
    7.663705e-06, 7.663699e-06, 7.663695e-06, 7.663692e-06, 7.663689e-06, 
    7.66368e-06, 7.663675e-06, 7.663665e-06, 7.663667e-06, 7.663663e-06, 
    7.663661e-06, 7.663655e-06, 7.663656e-06, 7.663654e-06, 7.663663e-06, 
    7.663657e-06, 7.663668e-06, 7.663665e-06, 7.663688e-06, 7.663697e-06, 
    7.663701e-06, 7.663704e-06, 7.663712e-06, 7.663706e-06, 7.663709e-06, 
    7.663703e-06, 7.6637e-06, 7.663702e-06, 7.663692e-06, 7.663696e-06, 
    7.663675e-06, 7.663684e-06, 7.663661e-06, 7.663666e-06, 7.66366e-06, 
    7.663663e-06, 7.663657e-06, 7.663662e-06, 7.663653e-06, 7.663652e-06, 
    7.663652e-06, 7.663647e-06, 7.663662e-06, 7.663657e-06, 7.663702e-06, 
    7.663702e-06, 7.663701e-06, 7.663706e-06, 7.663706e-06, 7.663712e-06, 
    7.663707e-06, 7.663705e-06, 7.6637e-06, 7.663697e-06, 7.663694e-06, 
    7.663689e-06, 7.663682e-06, 7.663672e-06, 7.663666e-06, 7.663662e-06, 
    7.663664e-06, 7.663662e-06, 7.663664e-06, 7.663666e-06, 7.663652e-06, 
    7.66366e-06, 7.663648e-06, 7.663649e-06, 7.663654e-06, 7.663649e-06, 
    7.663702e-06, 7.663703e-06, 7.663708e-06, 7.663704e-06, 7.663712e-06, 
    7.663707e-06, 7.663705e-06, 7.663695e-06, 7.663693e-06, 7.663692e-06, 
    7.663688e-06, 7.663683e-06, 7.663674e-06, 7.663667e-06, 7.663661e-06, 
    7.663661e-06, 7.663661e-06, 7.663659e-06, 7.663662e-06, 7.663659e-06, 
    7.663658e-06, 7.66366e-06, 7.663649e-06, 7.663652e-06, 7.663649e-06, 
    7.663651e-06, 7.663702e-06, 7.6637e-06, 7.663702e-06, 7.663699e-06, 
    7.663701e-06, 7.663692e-06, 7.66369e-06, 7.663678e-06, 7.663683e-06, 
    7.663675e-06, 7.663682e-06, 7.663682e-06, 7.663675e-06, 7.663682e-06, 
    7.663668e-06, 7.663677e-06, 7.663659e-06, 7.663669e-06, 7.663659e-06, 
    7.663661e-06, 7.663657e-06, 7.663654e-06, 7.663651e-06, 7.663644e-06, 
    7.663646e-06, 7.663641e-06, 7.663696e-06, 7.663692e-06, 7.663693e-06, 
    7.66369e-06, 7.663687e-06, 7.663682e-06, 7.663672e-06, 7.663676e-06, 
    7.66367e-06, 7.663668e-06, 7.663678e-06, 7.663672e-06, 7.663691e-06, 
    7.663687e-06, 7.663689e-06, 7.663696e-06, 7.663675e-06, 7.663685e-06, 
    7.663666e-06, 7.663672e-06, 7.663655e-06, 7.663663e-06, 7.663647e-06, 
    7.66364e-06, 7.663633e-06, 7.663625e-06, 7.663691e-06, 7.663693e-06, 
    7.663689e-06, 7.663683e-06, 7.663678e-06, 7.663672e-06, 7.663671e-06, 
    7.66367e-06, 7.663666e-06, 7.663663e-06, 7.663669e-06, 7.663662e-06, 
    7.663687e-06, 7.663674e-06, 7.663694e-06, 7.663688e-06, 7.663683e-06, 
    7.663685e-06, 7.663676e-06, 7.663674e-06, 7.663665e-06, 7.66367e-06, 
    7.663642e-06, 7.663654e-06, 7.66362e-06, 7.663629e-06, 7.663694e-06, 
    7.663691e-06, 7.663681e-06, 7.663685e-06, 7.663671e-06, 7.663667e-06, 
    7.663664e-06, 7.663661e-06, 7.663661e-06, 7.663658e-06, 7.663662e-06, 
    7.663658e-06, 7.663672e-06, 7.663665e-06, 7.663682e-06, 7.663678e-06, 
    7.66368e-06, 7.663682e-06, 7.663675e-06, 7.663669e-06, 7.663669e-06, 
    7.663667e-06, 7.663661e-06, 7.663671e-06, 7.66364e-06, 7.663659e-06, 
    7.663688e-06, 7.663682e-06, 7.663681e-06, 7.663683e-06, 7.663668e-06, 
    7.663673e-06, 7.663658e-06, 7.663662e-06, 7.663656e-06, 7.663659e-06, 
    7.66366e-06, 7.663663e-06, 7.663666e-06, 7.663673e-06, 7.663679e-06, 
    7.663682e-06, 7.663682e-06, 7.663677e-06, 7.663669e-06, 7.663661e-06, 
    7.663662e-06, 7.663656e-06, 7.663672e-06, 7.663665e-06, 7.663668e-06, 
    7.663662e-06, 7.663676e-06, 7.663663e-06, 7.663679e-06, 7.663678e-06, 
    7.663673e-06, 7.663665e-06, 7.663663e-06, 7.663661e-06, 7.663662e-06, 
    7.663668e-06, 7.663669e-06, 7.663673e-06, 7.663674e-06, 7.663678e-06, 
    7.663681e-06, 7.663678e-06, 7.663675e-06, 7.663668e-06, 7.663662e-06, 
    7.663654e-06, 7.663652e-06, 7.663644e-06, 7.663652e-06, 7.66364e-06, 
    7.66365e-06, 7.663632e-06, 7.663662e-06, 7.66365e-06, 7.663673e-06, 
    7.663671e-06, 7.663666e-06, 7.663655e-06, 7.663662e-06, 7.663654e-06, 
    7.663669e-06, 7.663677e-06, 7.663679e-06, 7.663682e-06, 7.663679e-06, 
    7.663679e-06, 7.663675e-06, 7.663677e-06, 7.663668e-06, 7.663672e-06, 
    7.66366e-06, 7.663654e-06, 7.663642e-06, 7.663632e-06, 7.663624e-06, 
    7.663621e-06, 7.66362e-06, 7.663619e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3_HR =
  5.325308e-14, 5.339687e-14, 5.336894e-14, 5.34848e-14, 5.342056e-14, 
    5.34964e-14, 5.328226e-14, 5.340256e-14, 5.332579e-14, 5.326606e-14, 
    5.370932e-14, 5.348997e-14, 5.393699e-14, 5.379734e-14, 5.41479e-14, 
    5.391524e-14, 5.419478e-14, 5.414124e-14, 5.430243e-14, 5.425628e-14, 
    5.446213e-14, 5.432373e-14, 5.456879e-14, 5.442912e-14, 5.445096e-14, 
    5.431915e-14, 5.353419e-14, 5.368202e-14, 5.352542e-14, 5.354651e-14, 
    5.353706e-14, 5.342187e-14, 5.336376e-14, 5.324212e-14, 5.326421e-14, 
    5.335357e-14, 5.3556e-14, 5.348735e-14, 5.366039e-14, 5.365648e-14, 
    5.384884e-14, 5.376214e-14, 5.408506e-14, 5.399339e-14, 5.425821e-14, 
    5.419164e-14, 5.425507e-14, 5.423584e-14, 5.425532e-14, 5.415769e-14, 
    5.419952e-14, 5.411359e-14, 5.377838e-14, 5.387698e-14, 5.358267e-14, 
    5.340533e-14, 5.328753e-14, 5.320385e-14, 5.321568e-14, 5.323823e-14, 
    5.335409e-14, 5.346298e-14, 5.35459e-14, 5.360133e-14, 5.365592e-14, 
    5.382092e-14, 5.390828e-14, 5.410357e-14, 5.406838e-14, 5.412801e-14, 
    5.418502e-14, 5.428062e-14, 5.426489e-14, 5.430698e-14, 5.412647e-14, 
    5.424645e-14, 5.404835e-14, 5.410254e-14, 5.36706e-14, 5.350588e-14, 
    5.343567e-14, 5.33743e-14, 5.322478e-14, 5.332804e-14, 5.328734e-14, 
    5.338419e-14, 5.344567e-14, 5.341527e-14, 5.360284e-14, 5.352994e-14, 
    5.391346e-14, 5.37484e-14, 5.417837e-14, 5.407561e-14, 5.4203e-14, 
    5.413802e-14, 5.424933e-14, 5.414915e-14, 5.432266e-14, 5.436039e-14, 
    5.43346e-14, 5.443368e-14, 5.414359e-14, 5.425506e-14, 5.341442e-14, 
    5.341937e-14, 5.344248e-14, 5.334086e-14, 5.333465e-14, 5.32415e-14, 
    5.33244e-14, 5.335968e-14, 5.344925e-14, 5.350217e-14, 5.355248e-14, 
    5.366301e-14, 5.378633e-14, 5.395862e-14, 5.408227e-14, 5.41651e-14, 
    5.411433e-14, 5.415915e-14, 5.410903e-14, 5.408554e-14, 5.434624e-14, 
    5.41999e-14, 5.441944e-14, 5.44073e-14, 5.430797e-14, 5.440867e-14, 
    5.342286e-14, 5.339432e-14, 5.329516e-14, 5.337277e-14, 5.323136e-14, 
    5.331051e-14, 5.335599e-14, 5.353143e-14, 5.356999e-14, 5.360568e-14, 
    5.367618e-14, 5.376658e-14, 5.392502e-14, 5.406271e-14, 5.418834e-14, 
    5.417914e-14, 5.418238e-14, 5.421041e-14, 5.414094e-14, 5.422182e-14, 
    5.423537e-14, 5.419991e-14, 5.440568e-14, 5.434693e-14, 5.440705e-14, 
    5.43688e-14, 5.34036e-14, 5.345161e-14, 5.342567e-14, 5.347445e-14, 
    5.344007e-14, 5.359281e-14, 5.363856e-14, 5.385252e-14, 5.376479e-14, 
    5.390443e-14, 5.3779e-14, 5.380122e-14, 5.390892e-14, 5.378579e-14, 
    5.405509e-14, 5.387252e-14, 5.42115e-14, 5.402933e-14, 5.422291e-14, 
    5.41878e-14, 5.424594e-14, 5.429798e-14, 5.436344e-14, 5.448409e-14, 
    5.445617e-14, 5.455704e-14, 5.352318e-14, 5.358538e-14, 5.357994e-14, 
    5.364503e-14, 5.369314e-14, 5.37974e-14, 5.396441e-14, 5.390164e-14, 
    5.401689e-14, 5.404e-14, 5.386492e-14, 5.397242e-14, 5.362702e-14, 
    5.368285e-14, 5.364964e-14, 5.352807e-14, 5.391607e-14, 5.371706e-14, 
    5.408431e-14, 5.397671e-14, 5.429055e-14, 5.413452e-14, 5.444079e-14, 
    5.457142e-14, 5.469439e-14, 5.483777e-14, 5.361935e-14, 5.357709e-14, 
    5.365277e-14, 5.375736e-14, 5.38544e-14, 5.398327e-14, 5.399646e-14, 
    5.402058e-14, 5.408304e-14, 5.413554e-14, 5.402818e-14, 5.41487e-14, 
    5.369574e-14, 5.393334e-14, 5.356109e-14, 5.367325e-14, 5.375121e-14, 
    5.371704e-14, 5.389447e-14, 5.393625e-14, 5.410582e-14, 5.401822e-14, 
    5.453916e-14, 5.430892e-14, 5.494694e-14, 5.476894e-14, 5.356232e-14, 
    5.361922e-14, 5.381702e-14, 5.372295e-14, 5.399188e-14, 5.405795e-14, 
    5.411169e-14, 5.418031e-14, 5.418774e-14, 5.422837e-14, 5.416177e-14, 
    5.422576e-14, 5.398354e-14, 5.409183e-14, 5.379446e-14, 5.386689e-14, 
    5.383359e-14, 5.379702e-14, 5.390983e-14, 5.402986e-14, 5.403247e-14, 
    5.40709e-14, 5.417911e-14, 5.399297e-14, 5.456876e-14, 5.421336e-14, 
    5.368124e-14, 5.379065e-14, 5.380633e-14, 5.376395e-14, 5.405136e-14, 
    5.394728e-14, 5.422739e-14, 5.415175e-14, 5.427568e-14, 5.42141e-14, 
    5.420504e-14, 5.412592e-14, 5.407663e-14, 5.395205e-14, 5.385059e-14, 
    5.377011e-14, 5.378882e-14, 5.387722e-14, 5.403721e-14, 5.418839e-14, 
    5.415527e-14, 5.426626e-14, 5.39724e-14, 5.409566e-14, 5.404803e-14, 
    5.417223e-14, 5.389996e-14, 5.41317e-14, 5.384064e-14, 5.38662e-14, 
    5.394522e-14, 5.410398e-14, 5.413916e-14, 5.417663e-14, 5.415352e-14, 
    5.404127e-14, 5.402289e-14, 5.394331e-14, 5.39213e-14, 5.386064e-14, 
    5.381036e-14, 5.385628e-14, 5.390448e-14, 5.404135e-14, 5.416451e-14, 
    5.429871e-14, 5.433155e-14, 5.448801e-14, 5.436059e-14, 5.457072e-14, 
    5.439199e-14, 5.470129e-14, 5.414519e-14, 5.438683e-14, 5.394883e-14, 
    5.39961e-14, 5.408147e-14, 5.427726e-14, 5.417165e-14, 5.429517e-14, 
    5.402218e-14, 5.388025e-14, 5.384356e-14, 5.377499e-14, 5.384513e-14, 
    5.383943e-14, 5.390651e-14, 5.388496e-14, 5.404589e-14, 5.395947e-14, 
    5.42048e-14, 5.429421e-14, 5.454645e-14, 5.470081e-14, 5.485782e-14, 
    5.492705e-14, 5.494812e-14, 5.495692e-14 ;

 LITTERC =
  5.976202e-05, 5.976187e-05, 5.97619e-05, 5.976178e-05, 5.976185e-05, 
    5.976177e-05, 5.976199e-05, 5.976186e-05, 5.976194e-05, 5.9762e-05, 
    5.976155e-05, 5.976178e-05, 5.976132e-05, 5.976146e-05, 5.976111e-05, 
    5.976134e-05, 5.976106e-05, 5.976111e-05, 5.976095e-05, 5.9761e-05, 
    5.976079e-05, 5.976093e-05, 5.976068e-05, 5.976082e-05, 5.97608e-05, 
    5.976094e-05, 5.976173e-05, 5.976158e-05, 5.976174e-05, 5.976172e-05, 
    5.976173e-05, 5.976185e-05, 5.97619e-05, 5.976203e-05, 5.976201e-05, 
    5.976191e-05, 5.976171e-05, 5.976178e-05, 5.97616e-05, 5.976161e-05, 
    5.976141e-05, 5.97615e-05, 5.976117e-05, 5.976126e-05, 5.9761e-05, 
    5.976106e-05, 5.9761e-05, 5.976102e-05, 5.9761e-05, 5.97611e-05, 
    5.976106e-05, 5.976114e-05, 5.976148e-05, 5.976138e-05, 5.976168e-05, 
    5.976186e-05, 5.976198e-05, 5.976206e-05, 5.976205e-05, 5.976203e-05, 
    5.976191e-05, 5.97618e-05, 5.976172e-05, 5.976166e-05, 5.976161e-05, 
    5.976144e-05, 5.976135e-05, 5.976115e-05, 5.976119e-05, 5.976113e-05, 
    5.976107e-05, 5.976097e-05, 5.976099e-05, 5.976095e-05, 5.976113e-05, 
    5.976101e-05, 5.976121e-05, 5.976115e-05, 5.976159e-05, 5.976176e-05, 
    5.976183e-05, 5.976189e-05, 5.976205e-05, 5.976194e-05, 5.976198e-05, 
    5.976188e-05, 5.976182e-05, 5.976185e-05, 5.976166e-05, 5.976174e-05, 
    5.976135e-05, 5.976151e-05, 5.976108e-05, 5.976118e-05, 5.976105e-05, 
    5.976112e-05, 5.976101e-05, 5.976111e-05, 5.976093e-05, 5.976089e-05, 
    5.976092e-05, 5.976082e-05, 5.976111e-05, 5.9761e-05, 5.976185e-05, 
    5.976185e-05, 5.976182e-05, 5.976193e-05, 5.976193e-05, 5.976203e-05, 
    5.976194e-05, 5.976191e-05, 5.976182e-05, 5.976176e-05, 5.976171e-05, 
    5.97616e-05, 5.976147e-05, 5.97613e-05, 5.976118e-05, 5.976109e-05, 
    5.976114e-05, 5.97611e-05, 5.976115e-05, 5.976117e-05, 5.976091e-05, 
    5.976106e-05, 5.976083e-05, 5.976085e-05, 5.976095e-05, 5.976085e-05, 
    5.976184e-05, 5.976187e-05, 5.976197e-05, 5.976189e-05, 5.976204e-05, 
    5.976196e-05, 5.976191e-05, 5.976173e-05, 5.976169e-05, 5.976166e-05, 
    5.976159e-05, 5.97615e-05, 5.976133e-05, 5.976119e-05, 5.976107e-05, 
    5.976108e-05, 5.976107e-05, 5.976105e-05, 5.976111e-05, 5.976103e-05, 
    5.976102e-05, 5.976106e-05, 5.976085e-05, 5.976091e-05, 5.976085e-05, 
    5.976089e-05, 5.976186e-05, 5.976181e-05, 5.976184e-05, 5.976179e-05, 
    5.976183e-05, 5.976167e-05, 5.976162e-05, 5.976141e-05, 5.97615e-05, 
    5.976135e-05, 5.976148e-05, 5.976146e-05, 5.976135e-05, 5.976147e-05, 
    5.97612e-05, 5.976139e-05, 5.976105e-05, 5.976123e-05, 5.976103e-05, 
    5.976107e-05, 5.976101e-05, 5.976096e-05, 5.976089e-05, 5.976077e-05, 
    5.97608e-05, 5.976069e-05, 5.976174e-05, 5.976168e-05, 5.976169e-05, 
    5.976162e-05, 5.976157e-05, 5.976146e-05, 5.976129e-05, 5.976136e-05, 
    5.976124e-05, 5.976122e-05, 5.976139e-05, 5.976129e-05, 5.976163e-05, 
    5.976158e-05, 5.976161e-05, 5.976174e-05, 5.976134e-05, 5.976154e-05, 
    5.976117e-05, 5.976128e-05, 5.976097e-05, 5.976112e-05, 5.976081e-05, 
    5.976068e-05, 5.976055e-05, 5.976041e-05, 5.976165e-05, 5.976169e-05, 
    5.976161e-05, 5.97615e-05, 5.976141e-05, 5.976127e-05, 5.976126e-05, 
    5.976124e-05, 5.976117e-05, 5.976112e-05, 5.976123e-05, 5.976111e-05, 
    5.976157e-05, 5.976133e-05, 5.97617e-05, 5.976159e-05, 5.976151e-05, 
    5.976154e-05, 5.976137e-05, 5.976132e-05, 5.976115e-05, 5.976124e-05, 
    5.976071e-05, 5.976095e-05, 5.97603e-05, 5.976048e-05, 5.97617e-05, 
    5.976165e-05, 5.976145e-05, 5.976154e-05, 5.976127e-05, 5.97612e-05, 
    5.976114e-05, 5.976107e-05, 5.976107e-05, 5.976103e-05, 5.97611e-05, 
    5.976103e-05, 5.976127e-05, 5.976117e-05, 5.976147e-05, 5.976139e-05, 
    5.976143e-05, 5.976146e-05, 5.976135e-05, 5.976123e-05, 5.976123e-05, 
    5.976119e-05, 5.976108e-05, 5.976127e-05, 5.976068e-05, 5.976104e-05, 
    5.976158e-05, 5.976147e-05, 5.976146e-05, 5.97615e-05, 5.976121e-05, 
    5.976131e-05, 5.976103e-05, 5.97611e-05, 5.976098e-05, 5.976104e-05, 
    5.976105e-05, 5.976113e-05, 5.976118e-05, 5.976131e-05, 5.976141e-05, 
    5.976149e-05, 5.976147e-05, 5.976138e-05, 5.976122e-05, 5.976107e-05, 
    5.97611e-05, 5.976099e-05, 5.976129e-05, 5.976116e-05, 5.976121e-05, 
    5.976109e-05, 5.976136e-05, 5.976113e-05, 5.976142e-05, 5.976139e-05, 
    5.976131e-05, 5.976115e-05, 5.976112e-05, 5.976108e-05, 5.97611e-05, 
    5.976122e-05, 5.976123e-05, 5.976131e-05, 5.976134e-05, 5.97614e-05, 
    5.976145e-05, 5.976141e-05, 5.976135e-05, 5.976122e-05, 5.976109e-05, 
    5.976095e-05, 5.976092e-05, 5.976076e-05, 5.976089e-05, 5.976068e-05, 
    5.976086e-05, 5.976055e-05, 5.976111e-05, 5.976087e-05, 5.976131e-05, 
    5.976126e-05, 5.976118e-05, 5.976098e-05, 5.976109e-05, 5.976096e-05, 
    5.976123e-05, 5.976138e-05, 5.976142e-05, 5.976149e-05, 5.976142e-05, 
    5.976142e-05, 5.976135e-05, 5.976138e-05, 5.976121e-05, 5.97613e-05, 
    5.976105e-05, 5.976096e-05, 5.97607e-05, 5.976055e-05, 5.976039e-05, 
    5.976032e-05, 5.97603e-05, 5.976029e-05 ;

 LITTERC_HR =
  8.591897e-13, 8.615078e-13, 8.610575e-13, 8.629254e-13, 8.618897e-13, 
    8.631123e-13, 8.596602e-13, 8.615995e-13, 8.603619e-13, 8.593989e-13, 
    8.66545e-13, 8.630088e-13, 8.702151e-13, 8.679639e-13, 8.736153e-13, 
    8.698645e-13, 8.743711e-13, 8.73508e-13, 8.761065e-13, 8.753624e-13, 
    8.78681e-13, 8.764498e-13, 8.804005e-13, 8.781488e-13, 8.785009e-13, 
    8.76376e-13, 8.637216e-13, 8.661048e-13, 8.635801e-13, 8.639202e-13, 
    8.637678e-13, 8.619109e-13, 8.60974e-13, 8.590129e-13, 8.593692e-13, 
    8.608098e-13, 8.640731e-13, 8.629664e-13, 8.65756e-13, 8.656931e-13, 
    8.687941e-13, 8.673965e-13, 8.726022e-13, 8.711244e-13, 8.753935e-13, 
    8.743204e-13, 8.75343e-13, 8.750331e-13, 8.75347e-13, 8.737731e-13, 
    8.744475e-13, 8.730623e-13, 8.676582e-13, 8.692477e-13, 8.645031e-13, 
    8.616442e-13, 8.597452e-13, 8.58396e-13, 8.585868e-13, 8.589503e-13, 
    8.608182e-13, 8.625737e-13, 8.639103e-13, 8.648039e-13, 8.65684e-13, 
    8.683441e-13, 8.697523e-13, 8.729006e-13, 8.723333e-13, 8.732947e-13, 
    8.742137e-13, 8.757548e-13, 8.755013e-13, 8.761798e-13, 8.732698e-13, 
    8.75204e-13, 8.720105e-13, 8.72884e-13, 8.659207e-13, 8.632651e-13, 
    8.621332e-13, 8.611439e-13, 8.587334e-13, 8.603982e-13, 8.59742e-13, 
    8.613034e-13, 8.622946e-13, 8.618045e-13, 8.648283e-13, 8.636531e-13, 
    8.698358e-13, 8.671749e-13, 8.741065e-13, 8.724498e-13, 8.745035e-13, 
    8.734559e-13, 8.752503e-13, 8.736355e-13, 8.764325e-13, 8.770408e-13, 
    8.766251e-13, 8.782224e-13, 8.735458e-13, 8.753427e-13, 8.617907e-13, 
    8.618706e-13, 8.622432e-13, 8.606048e-13, 8.605048e-13, 8.59003e-13, 
    8.603395e-13, 8.609082e-13, 8.623522e-13, 8.632054e-13, 8.640164e-13, 
    8.657984e-13, 8.677864e-13, 8.70564e-13, 8.725572e-13, 8.738925e-13, 
    8.73074e-13, 8.737966e-13, 8.729887e-13, 8.7261e-13, 8.768127e-13, 
    8.744536e-13, 8.779927e-13, 8.777971e-13, 8.761959e-13, 8.778192e-13, 
    8.619267e-13, 8.614667e-13, 8.598681e-13, 8.611193e-13, 8.588395e-13, 
    8.601155e-13, 8.608488e-13, 8.636771e-13, 8.642987e-13, 8.648741e-13, 
    8.660107e-13, 8.67468e-13, 8.700222e-13, 8.72242e-13, 8.742672e-13, 
    8.74119e-13, 8.741711e-13, 8.746231e-13, 8.735031e-13, 8.748069e-13, 
    8.750254e-13, 8.744537e-13, 8.777709e-13, 8.768238e-13, 8.77793e-13, 
    8.771764e-13, 8.616163e-13, 8.623903e-13, 8.619721e-13, 8.627584e-13, 
    8.622043e-13, 8.646666e-13, 8.654043e-13, 8.688535e-13, 8.674392e-13, 
    8.696903e-13, 8.676682e-13, 8.680265e-13, 8.697626e-13, 8.677777e-13, 
    8.721191e-13, 8.691759e-13, 8.746406e-13, 8.717039e-13, 8.748245e-13, 
    8.742585e-13, 8.751958e-13, 8.760347e-13, 8.7709e-13, 8.79035e-13, 
    8.785849e-13, 8.802109e-13, 8.63544e-13, 8.645469e-13, 8.644591e-13, 
    8.655085e-13, 8.66284e-13, 8.679648e-13, 8.706572e-13, 8.696453e-13, 
    8.715032e-13, 8.718759e-13, 8.690534e-13, 8.707863e-13, 8.652181e-13, 
    8.661182e-13, 8.655827e-13, 8.636229e-13, 8.698778e-13, 8.666697e-13, 
    8.725901e-13, 8.708555e-13, 8.75915e-13, 8.733995e-13, 8.783369e-13, 
    8.804428e-13, 8.824252e-13, 8.847366e-13, 8.650945e-13, 8.644133e-13, 
    8.656333e-13, 8.673193e-13, 8.688838e-13, 8.709612e-13, 8.71174e-13, 
    8.715628e-13, 8.725696e-13, 8.73416e-13, 8.716852e-13, 8.736282e-13, 
    8.663259e-13, 8.701563e-13, 8.641552e-13, 8.659634e-13, 8.672201e-13, 
    8.666694e-13, 8.695298e-13, 8.702032e-13, 8.729369e-13, 8.715247e-13, 
    8.799228e-13, 8.762111e-13, 8.864965e-13, 8.83627e-13, 8.641751e-13, 
    8.650924e-13, 8.682811e-13, 8.667646e-13, 8.711001e-13, 8.721653e-13, 
    8.730316e-13, 8.741377e-13, 8.742575e-13, 8.749126e-13, 8.738389e-13, 
    8.748704e-13, 8.709657e-13, 8.727113e-13, 8.679175e-13, 8.690851e-13, 
    8.685482e-13, 8.679588e-13, 8.697773e-13, 8.717123e-13, 8.717544e-13, 
    8.723739e-13, 8.741185e-13, 8.711177e-13, 8.803999e-13, 8.746705e-13, 
    8.660921e-13, 8.67856e-13, 8.681088e-13, 8.674256e-13, 8.720589e-13, 
    8.703811e-13, 8.748967e-13, 8.736773e-13, 8.756752e-13, 8.746825e-13, 
    8.745364e-13, 8.73261e-13, 8.724663e-13, 8.704579e-13, 8.688223e-13, 
    8.675248e-13, 8.678266e-13, 8.692517e-13, 8.718308e-13, 8.742679e-13, 
    8.737341e-13, 8.755234e-13, 8.70786e-13, 8.727731e-13, 8.720053e-13, 
    8.740076e-13, 8.696182e-13, 8.733541e-13, 8.686619e-13, 8.690739e-13, 
    8.703478e-13, 8.729073e-13, 8.734744e-13, 8.740784e-13, 8.737059e-13, 
    8.718964e-13, 8.716001e-13, 8.703171e-13, 8.699623e-13, 8.689842e-13, 
    8.681739e-13, 8.689141e-13, 8.696911e-13, 8.718975e-13, 8.73883e-13, 
    8.760465e-13, 8.765759e-13, 8.790982e-13, 8.77044e-13, 8.804316e-13, 
    8.775502e-13, 8.825364e-13, 8.735716e-13, 8.77467e-13, 8.70406e-13, 
    8.711681e-13, 8.725444e-13, 8.757007e-13, 8.739981e-13, 8.759895e-13, 
    8.715886e-13, 8.693005e-13, 8.68709e-13, 8.676036e-13, 8.687343e-13, 
    8.686424e-13, 8.697238e-13, 8.693764e-13, 8.719707e-13, 8.705776e-13, 
    8.745325e-13, 8.75974e-13, 8.800403e-13, 8.825286e-13, 8.850598e-13, 
    8.861758e-13, 8.865154e-13, 8.866573e-13 ;

 LITTERC_LOSS =
  1.59121e-12, 1.595503e-12, 1.594669e-12, 1.598129e-12, 1.596211e-12, 
    1.598475e-12, 1.592082e-12, 1.595673e-12, 1.593381e-12, 1.591598e-12, 
    1.604832e-12, 1.598283e-12, 1.61163e-12, 1.60746e-12, 1.617927e-12, 
    1.61098e-12, 1.619326e-12, 1.617728e-12, 1.62254e-12, 1.621162e-12, 
    1.627308e-12, 1.623176e-12, 1.630493e-12, 1.626323e-12, 1.626975e-12, 
    1.62304e-12, 1.599603e-12, 1.604017e-12, 1.599341e-12, 1.599971e-12, 
    1.599689e-12, 1.59625e-12, 1.594515e-12, 1.590883e-12, 1.591543e-12, 
    1.594211e-12, 1.600254e-12, 1.598205e-12, 1.603371e-12, 1.603255e-12, 
    1.608998e-12, 1.606409e-12, 1.61605e-12, 1.613314e-12, 1.62122e-12, 
    1.619233e-12, 1.621126e-12, 1.620552e-12, 1.621134e-12, 1.618219e-12, 
    1.619468e-12, 1.616902e-12, 1.606894e-12, 1.609838e-12, 1.601051e-12, 
    1.595756e-12, 1.592239e-12, 1.58974e-12, 1.590094e-12, 1.590767e-12, 
    1.594226e-12, 1.597477e-12, 1.599953e-12, 1.601608e-12, 1.603238e-12, 
    1.608164e-12, 1.610772e-12, 1.616603e-12, 1.615552e-12, 1.617333e-12, 
    1.619035e-12, 1.621889e-12, 1.62142e-12, 1.622676e-12, 1.617287e-12, 
    1.620869e-12, 1.614954e-12, 1.616572e-12, 1.603676e-12, 1.598758e-12, 
    1.596662e-12, 1.59483e-12, 1.590365e-12, 1.593448e-12, 1.592233e-12, 
    1.595125e-12, 1.596961e-12, 1.596053e-12, 1.601653e-12, 1.599477e-12, 
    1.610927e-12, 1.605999e-12, 1.618836e-12, 1.615768e-12, 1.619572e-12, 
    1.617631e-12, 1.620955e-12, 1.617964e-12, 1.623144e-12, 1.624271e-12, 
    1.623501e-12, 1.626459e-12, 1.617798e-12, 1.621126e-12, 1.596027e-12, 
    1.596175e-12, 1.596865e-12, 1.593831e-12, 1.593646e-12, 1.590864e-12, 
    1.59334e-12, 1.594393e-12, 1.597067e-12, 1.598647e-12, 1.600149e-12, 
    1.60345e-12, 1.607131e-12, 1.612276e-12, 1.615967e-12, 1.61844e-12, 
    1.616924e-12, 1.618262e-12, 1.616766e-12, 1.616065e-12, 1.623848e-12, 
    1.619479e-12, 1.626034e-12, 1.625671e-12, 1.622706e-12, 1.625712e-12, 
    1.596279e-12, 1.595427e-12, 1.592467e-12, 1.594784e-12, 1.590562e-12, 
    1.592925e-12, 1.594283e-12, 1.599521e-12, 1.600672e-12, 1.601738e-12, 
    1.603843e-12, 1.606542e-12, 1.611272e-12, 1.615383e-12, 1.619134e-12, 
    1.618859e-12, 1.618956e-12, 1.619793e-12, 1.617719e-12, 1.620133e-12, 
    1.620538e-12, 1.619479e-12, 1.625623e-12, 1.623869e-12, 1.625664e-12, 
    1.624522e-12, 1.595704e-12, 1.597138e-12, 1.596363e-12, 1.59782e-12, 
    1.596793e-12, 1.601353e-12, 1.60272e-12, 1.609108e-12, 1.606488e-12, 
    1.610658e-12, 1.606913e-12, 1.607576e-12, 1.610791e-12, 1.607115e-12, 
    1.615156e-12, 1.609705e-12, 1.619826e-12, 1.614387e-12, 1.620166e-12, 
    1.619118e-12, 1.620854e-12, 1.622407e-12, 1.624362e-12, 1.627964e-12, 
    1.62713e-12, 1.630142e-12, 1.599275e-12, 1.601132e-12, 1.600969e-12, 
    1.602913e-12, 1.604349e-12, 1.607462e-12, 1.612448e-12, 1.610574e-12, 
    1.614015e-12, 1.614705e-12, 1.609478e-12, 1.612687e-12, 1.602375e-12, 
    1.604042e-12, 1.60305e-12, 1.599421e-12, 1.611005e-12, 1.605063e-12, 
    1.616028e-12, 1.612815e-12, 1.622186e-12, 1.617527e-12, 1.626671e-12, 
    1.630571e-12, 1.634243e-12, 1.638524e-12, 1.602146e-12, 1.600884e-12, 
    1.603144e-12, 1.606266e-12, 1.609164e-12, 1.613011e-12, 1.613405e-12, 
    1.614125e-12, 1.61599e-12, 1.617558e-12, 1.614352e-12, 1.61795e-12, 
    1.604427e-12, 1.611521e-12, 1.600406e-12, 1.603755e-12, 1.606083e-12, 
    1.605063e-12, 1.61036e-12, 1.611607e-12, 1.61667e-12, 1.614055e-12, 
    1.629608e-12, 1.622734e-12, 1.641783e-12, 1.636469e-12, 1.600443e-12, 
    1.602142e-12, 1.608048e-12, 1.605239e-12, 1.613269e-12, 1.615241e-12, 
    1.616846e-12, 1.618894e-12, 1.619116e-12, 1.620329e-12, 1.618341e-12, 
    1.620251e-12, 1.61302e-12, 1.616252e-12, 1.607374e-12, 1.609537e-12, 
    1.608542e-12, 1.607451e-12, 1.610819e-12, 1.614402e-12, 1.61448e-12, 
    1.615628e-12, 1.618859e-12, 1.613301e-12, 1.630492e-12, 1.619881e-12, 
    1.603994e-12, 1.60726e-12, 1.607728e-12, 1.606463e-12, 1.615044e-12, 
    1.611937e-12, 1.6203e-12, 1.618042e-12, 1.621742e-12, 1.619903e-12, 
    1.619633e-12, 1.617271e-12, 1.615799e-12, 1.612079e-12, 1.60905e-12, 
    1.606647e-12, 1.607206e-12, 1.609845e-12, 1.614622e-12, 1.619135e-12, 
    1.618147e-12, 1.621461e-12, 1.612687e-12, 1.616367e-12, 1.614945e-12, 
    1.618653e-12, 1.610524e-12, 1.617443e-12, 1.608753e-12, 1.609516e-12, 
    1.611875e-12, 1.616615e-12, 1.617666e-12, 1.618784e-12, 1.618094e-12, 
    1.614743e-12, 1.614194e-12, 1.611818e-12, 1.611161e-12, 1.60935e-12, 
    1.607849e-12, 1.60922e-12, 1.610659e-12, 1.614745e-12, 1.618422e-12, 
    1.622429e-12, 1.62341e-12, 1.628081e-12, 1.624277e-12, 1.630551e-12, 
    1.625214e-12, 1.634449e-12, 1.617846e-12, 1.62506e-12, 1.611983e-12, 
    1.613394e-12, 1.615943e-12, 1.621789e-12, 1.618636e-12, 1.622324e-12, 
    1.614173e-12, 1.609935e-12, 1.60884e-12, 1.606793e-12, 1.608887e-12, 
    1.608717e-12, 1.61072e-12, 1.610076e-12, 1.614881e-12, 1.612301e-12, 
    1.619625e-12, 1.622295e-12, 1.629826e-12, 1.634434e-12, 1.639122e-12, 
    1.641189e-12, 1.641818e-12, 1.642081e-12 ;

 LIVECROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVECROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 MEG_acetaldehyde =
  3.91629e-18, 3.914856e-18, 3.915128e-18, 3.913988e-18, 3.91461e-18, 
    3.913872e-18, 3.915987e-18, 3.914811e-18, 3.915554e-18, 3.916144e-18, 
    3.911814e-18, 3.913934e-18, 3.909504e-18, 3.91087e-18, 3.907407e-18, 
    3.909732e-18, 3.906934e-18, 3.907446e-18, 3.905838e-18, 3.906296e-18, 
    3.904299e-18, 3.905625e-18, 3.903221e-18, 3.904601e-18, 3.904395e-18, 
    3.905673e-18, 3.913481e-18, 3.912087e-18, 3.91357e-18, 3.91337e-18, 
    3.913454e-18, 3.914607e-18, 3.915207e-18, 3.916381e-18, 3.916163e-18, 
    3.91529e-18, 3.913279e-18, 3.913943e-18, 3.912217e-18, 3.912255e-18, 
    3.910356e-18, 3.911212e-18, 3.908005e-18, 3.908909e-18, 3.906277e-18, 
    3.906942e-18, 3.906313e-18, 3.9065e-18, 3.90631e-18, 3.907284e-18, 
    3.906869e-18, 3.907718e-18, 3.911057e-18, 3.910083e-18, 3.913006e-18, 
    3.914808e-18, 3.91594e-18, 3.916765e-18, 3.916649e-18, 3.916432e-18, 
    3.915285e-18, 3.914186e-18, 3.913357e-18, 3.912807e-18, 3.912261e-18, 
    3.910683e-18, 3.909789e-18, 3.907836e-18, 3.908165e-18, 3.90759e-18, 
    3.907007e-18, 3.906062e-18, 3.906214e-18, 3.905803e-18, 3.907588e-18, 
    3.90641e-18, 3.908358e-18, 3.907827e-18, 3.912205e-18, 3.913759e-18, 
    3.9145e-18, 3.915079e-18, 3.91656e-18, 3.915543e-18, 3.915946e-18, 
    3.914967e-18, 3.914359e-18, 3.914656e-18, 3.912791e-18, 3.913519e-18, 
    3.909737e-18, 3.911363e-18, 3.907075e-18, 3.908095e-18, 3.906827e-18, 
    3.90747e-18, 3.906377e-18, 3.90736e-18, 3.905643e-18, 3.90528e-18, 
    3.90553e-18, 3.904539e-18, 3.907417e-18, 3.906322e-18, 3.914668e-18, 
    3.914621e-18, 3.914387e-18, 3.915417e-18, 3.915475e-18, 3.916392e-18, 
    3.915567e-18, 3.915224e-18, 3.914316e-18, 3.913797e-18, 3.913298e-18, 
    3.9122e-18, 3.91099e-18, 3.909275e-18, 3.90803e-18, 3.907201e-18, 
    3.907703e-18, 3.907261e-18, 3.907759e-18, 3.907989e-18, 3.905422e-18, 
    3.90687e-18, 3.904682e-18, 3.904799e-18, 3.905797e-18, 3.904786e-18, 
    3.914586e-18, 3.914864e-18, 3.915861e-18, 3.915081e-18, 3.91649e-18, 
    3.915713e-18, 3.915272e-18, 3.913524e-18, 3.913119e-18, 3.912771e-18, 
    3.912064e-18, 3.911169e-18, 3.909606e-18, 3.908234e-18, 3.90697e-18, 
    3.907061e-18, 3.907029e-18, 3.906757e-18, 3.907444e-18, 3.906643e-18, 
    3.906517e-18, 3.90686e-18, 3.904816e-18, 3.905398e-18, 3.904802e-18, 
    3.905178e-18, 3.914771e-18, 3.914298e-18, 3.914555e-18, 3.914078e-18, 
    3.914421e-18, 3.912919e-18, 3.91247e-18, 3.910342e-18, 3.911192e-18, 
    3.909815e-18, 3.911044e-18, 3.910832e-18, 3.909809e-18, 3.910972e-18, 
    3.908327e-18, 3.910153e-18, 3.906746e-18, 3.908604e-18, 3.906632e-18, 
    3.906975e-18, 3.906397e-18, 3.90589e-18, 3.905235e-18, 3.904056e-18, 
    3.904325e-18, 3.903324e-18, 3.913585e-18, 3.912982e-18, 3.913018e-18, 
    3.912374e-18, 3.911902e-18, 3.910858e-18, 3.909207e-18, 3.909822e-18, 
    3.908674e-18, 3.90845e-18, 3.910184e-18, 3.909135e-18, 3.912564e-18, 
    3.912028e-18, 3.912335e-18, 3.913548e-18, 3.909704e-18, 3.911685e-18, 
    3.908013e-18, 3.909081e-18, 3.905965e-18, 3.90753e-18, 3.904477e-18, 
    3.90322e-18, 3.901958e-18, 3.900578e-18, 3.912633e-18, 3.913045e-18, 
    3.912292e-18, 3.911283e-18, 3.910299e-18, 3.909019e-18, 3.908878e-18, 
    3.908644e-18, 3.908015e-18, 3.907496e-18, 3.908586e-18, 3.907364e-18, 
    3.911938e-18, 3.909524e-18, 3.913217e-18, 3.912127e-18, 3.911335e-18, 
    3.911665e-18, 3.909888e-18, 3.909476e-18, 3.907808e-18, 3.90866e-18, 
    3.903545e-18, 3.905807e-18, 3.899472e-18, 3.901249e-18, 3.913194e-18, 
    3.912627e-18, 3.910681e-18, 3.911604e-18, 3.908924e-18, 3.908273e-18, 
    3.907729e-18, 3.907063e-18, 3.906978e-18, 3.906582e-18, 3.907234e-18, 
    3.906601e-18, 3.909016e-18, 3.907933e-18, 3.910883e-18, 3.910174e-18, 
    3.910494e-18, 3.910858e-18, 3.909737e-18, 3.908574e-18, 3.908521e-18, 
    3.908153e-18, 3.907165e-18, 3.908912e-18, 3.903304e-18, 3.906811e-18, 
    3.91201e-18, 3.910958e-18, 3.910774e-18, 3.911187e-18, 3.90834e-18, 
    3.909374e-18, 3.906588e-18, 3.907334e-18, 3.906104e-18, 3.906717e-18, 
    3.906809e-18, 3.907591e-18, 3.908086e-18, 3.909332e-18, 3.910339e-18, 
    3.911124e-18, 3.910939e-18, 3.910077e-18, 3.908496e-18, 3.906984e-18, 
    3.907318e-18, 3.906197e-18, 3.909119e-18, 3.907907e-18, 3.908385e-18, 
    3.907135e-18, 3.909844e-18, 3.907621e-18, 3.910424e-18, 3.910172e-18, 
    3.909394e-18, 3.907844e-18, 3.907459e-18, 3.9071e-18, 3.907316e-18, 
    3.908451e-18, 3.908624e-18, 3.909407e-18, 3.909636e-18, 3.910224e-18, 
    3.910725e-18, 3.910275e-18, 3.909808e-18, 3.908439e-18, 3.907222e-18, 
    3.905887e-18, 3.90555e-18, 3.904063e-18, 3.905311e-18, 3.90329e-18, 
    3.905065e-18, 3.901966e-18, 3.907451e-18, 3.905062e-18, 3.909349e-18, 
    3.90888e-18, 3.908061e-18, 3.906126e-18, 3.90714e-18, 3.90594e-18, 
    3.908629e-18, 3.91006e-18, 3.910397e-18, 3.911081e-18, 3.910381e-18, 
    3.910437e-18, 3.909769e-18, 3.909982e-18, 3.908393e-18, 3.909245e-18, 
    3.906819e-18, 3.905943e-18, 3.903439e-18, 3.901925e-18, 3.900341e-18, 
    3.899658e-18, 3.899448e-18, 3.899361e-18 ;

 MEG_acetic_acid =
  5.874435e-19, 5.872284e-19, 5.872692e-19, 5.870982e-19, 5.871915e-19, 
    5.870807e-19, 5.87398e-19, 5.872215e-19, 5.873331e-19, 5.874216e-19, 
    5.867721e-19, 5.8709e-19, 5.864256e-19, 5.866305e-19, 5.86111e-19, 
    5.864598e-19, 5.8604e-19, 5.861169e-19, 5.858756e-19, 5.859445e-19, 
    5.856448e-19, 5.858438e-19, 5.854832e-19, 5.856901e-19, 5.856593e-19, 
    5.85851e-19, 5.870221e-19, 5.86813e-19, 5.870354e-19, 5.870054e-19, 
    5.87018e-19, 5.87191e-19, 5.87281e-19, 5.874571e-19, 5.874244e-19, 
    5.872935e-19, 5.869918e-19, 5.870914e-19, 5.868325e-19, 5.868383e-19, 
    5.865534e-19, 5.866818e-19, 5.862008e-19, 5.863364e-19, 5.859415e-19, 
    5.860413e-19, 5.859469e-19, 5.85975e-19, 5.859465e-19, 5.860927e-19, 
    5.860303e-19, 5.861577e-19, 5.866585e-19, 5.865125e-19, 5.869508e-19, 
    5.872212e-19, 5.87391e-19, 5.875147e-19, 5.874973e-19, 5.874648e-19, 
    5.872928e-19, 5.871278e-19, 5.870034e-19, 5.86921e-19, 5.868391e-19, 
    5.866024e-19, 5.864683e-19, 5.861753e-19, 5.862247e-19, 5.861384e-19, 
    5.860511e-19, 5.859092e-19, 5.85932e-19, 5.858704e-19, 5.861381e-19, 
    5.859614e-19, 5.862537e-19, 5.861741e-19, 5.868308e-19, 5.870639e-19, 
    5.87175e-19, 5.872619e-19, 5.874841e-19, 5.873314e-19, 5.873919e-19, 
    5.872451e-19, 5.871538e-19, 5.871984e-19, 5.869187e-19, 5.870279e-19, 
    5.864605e-19, 5.867044e-19, 5.860612e-19, 5.862143e-19, 5.860241e-19, 
    5.861204e-19, 5.859565e-19, 5.861039e-19, 5.858464e-19, 5.857919e-19, 
    5.858294e-19, 5.856808e-19, 5.861125e-19, 5.859482e-19, 5.872003e-19, 
    5.871931e-19, 5.871581e-19, 5.873125e-19, 5.873212e-19, 5.874587e-19, 
    5.87335e-19, 5.872836e-19, 5.871474e-19, 5.870696e-19, 5.869947e-19, 
    5.8683e-19, 5.866485e-19, 5.863913e-19, 5.862045e-19, 5.860802e-19, 
    5.861555e-19, 5.860891e-19, 5.861639e-19, 5.861983e-19, 5.858132e-19, 
    5.860305e-19, 5.857022e-19, 5.857199e-19, 5.858695e-19, 5.857179e-19, 
    5.871878e-19, 5.872296e-19, 5.873791e-19, 5.87262e-19, 5.874735e-19, 
    5.873569e-19, 5.872908e-19, 5.870286e-19, 5.869677e-19, 5.869157e-19, 
    5.868096e-19, 5.866753e-19, 5.864409e-19, 5.86235e-19, 5.860454e-19, 
    5.860591e-19, 5.860544e-19, 5.860135e-19, 5.861167e-19, 5.859964e-19, 
    5.859775e-19, 5.860289e-19, 5.857224e-19, 5.858097e-19, 5.857203e-19, 
    5.857767e-19, 5.872156e-19, 5.871447e-19, 5.871833e-19, 5.871116e-19, 
    5.871631e-19, 5.869379e-19, 5.868704e-19, 5.865513e-19, 5.866787e-19, 
    5.864722e-19, 5.866567e-19, 5.866247e-19, 5.864713e-19, 5.866457e-19, 
    5.86249e-19, 5.86523e-19, 5.860119e-19, 5.862905e-19, 5.859948e-19, 
    5.860462e-19, 5.859596e-19, 5.858835e-19, 5.857853e-19, 5.856083e-19, 
    5.856487e-19, 5.854986e-19, 5.870378e-19, 5.869473e-19, 5.869526e-19, 
    5.868561e-19, 5.867853e-19, 5.866287e-19, 5.86381e-19, 5.864733e-19, 
    5.863011e-19, 5.862675e-19, 5.865275e-19, 5.863703e-19, 5.868846e-19, 
    5.868041e-19, 5.868502e-19, 5.870321e-19, 5.864556e-19, 5.867528e-19, 
    5.862019e-19, 5.863621e-19, 5.858947e-19, 5.861295e-19, 5.856715e-19, 
    5.854829e-19, 5.852937e-19, 5.850867e-19, 5.86895e-19, 5.869568e-19, 
    5.868438e-19, 5.866925e-19, 5.865448e-19, 5.863528e-19, 5.863317e-19, 
    5.862966e-19, 5.862022e-19, 5.861243e-19, 5.862879e-19, 5.861046e-19, 
    5.867906e-19, 5.864287e-19, 5.869826e-19, 5.86819e-19, 5.867002e-19, 
    5.867497e-19, 5.864832e-19, 5.864214e-19, 5.861713e-19, 5.86299e-19, 
    5.855317e-19, 5.85871e-19, 5.849208e-19, 5.851874e-19, 5.86979e-19, 
    5.86894e-19, 5.866022e-19, 5.867405e-19, 5.863386e-19, 5.862409e-19, 
    5.861594e-19, 5.860595e-19, 5.860468e-19, 5.859873e-19, 5.860851e-19, 
    5.859902e-19, 5.863524e-19, 5.8619e-19, 5.866324e-19, 5.865261e-19, 
    5.865741e-19, 5.866287e-19, 5.864606e-19, 5.86286e-19, 5.862781e-19, 
    5.862228e-19, 5.860747e-19, 5.863368e-19, 5.854956e-19, 5.860216e-19, 
    5.868016e-19, 5.866437e-19, 5.866161e-19, 5.866781e-19, 5.862509e-19, 
    5.864061e-19, 5.859881e-19, 5.861001e-19, 5.859157e-19, 5.860076e-19, 
    5.860213e-19, 5.861386e-19, 5.862128e-19, 5.863998e-19, 5.865508e-19, 
    5.866686e-19, 5.866409e-19, 5.865114e-19, 5.862743e-19, 5.860475e-19, 
    5.860977e-19, 5.859296e-19, 5.863678e-19, 5.86186e-19, 5.862576e-19, 
    5.860703e-19, 5.864766e-19, 5.861431e-19, 5.865635e-19, 5.865257e-19, 
    5.864091e-19, 5.861765e-19, 5.861189e-19, 5.86065e-19, 5.860974e-19, 
    5.862676e-19, 5.862936e-19, 5.864109e-19, 5.864454e-19, 5.865336e-19, 
    5.866087e-19, 5.865412e-19, 5.864711e-19, 5.862658e-19, 5.860832e-19, 
    5.858831e-19, 5.858325e-19, 5.856094e-19, 5.857966e-19, 5.854934e-19, 
    5.857597e-19, 5.852948e-19, 5.861176e-19, 5.857593e-19, 5.864024e-19, 
    5.86332e-19, 5.86209e-19, 5.859189e-19, 5.860711e-19, 5.85891e-19, 
    5.862943e-19, 5.865091e-19, 5.865595e-19, 5.866622e-19, 5.865571e-19, 
    5.865655e-19, 5.864653e-19, 5.864973e-19, 5.862589e-19, 5.863867e-19, 
    5.860228e-19, 5.858914e-19, 5.855158e-19, 5.852887e-19, 5.850512e-19, 
    5.849487e-19, 5.849171e-19, 5.849041e-19 ;

 MEG_acetone =
  1.22078e-16, 1.220548e-16, 1.220592e-16, 1.220408e-16, 1.220509e-16, 
    1.220389e-16, 1.220731e-16, 1.220541e-16, 1.220661e-16, 1.220757e-16, 
    1.220056e-16, 1.220399e-16, 1.219683e-16, 1.219904e-16, 1.219344e-16, 
    1.21972e-16, 1.219267e-16, 1.21935e-16, 1.21909e-16, 1.219164e-16, 
    1.218842e-16, 1.219056e-16, 1.218668e-16, 1.218891e-16, 1.218858e-16, 
    1.219064e-16, 1.220326e-16, 1.2201e-16, 1.22034e-16, 1.220308e-16, 
    1.220321e-16, 1.220508e-16, 1.220605e-16, 1.220795e-16, 1.22076e-16, 
    1.220619e-16, 1.220293e-16, 1.220401e-16, 1.220121e-16, 1.220128e-16, 
    1.21982e-16, 1.219959e-16, 1.21944e-16, 1.219587e-16, 1.219161e-16, 
    1.219269e-16, 1.219167e-16, 1.219197e-16, 1.219167e-16, 1.219324e-16, 
    1.219257e-16, 1.219394e-16, 1.219934e-16, 1.219776e-16, 1.220249e-16, 
    1.22054e-16, 1.220724e-16, 1.220857e-16, 1.220838e-16, 1.220803e-16, 
    1.220618e-16, 1.22044e-16, 1.220306e-16, 1.220217e-16, 1.220129e-16, 
    1.219873e-16, 1.219729e-16, 1.219413e-16, 1.219466e-16, 1.219373e-16, 
    1.219279e-16, 1.219126e-16, 1.219151e-16, 1.219085e-16, 1.219373e-16, 
    1.219183e-16, 1.219498e-16, 1.219412e-16, 1.220119e-16, 1.220371e-16, 
    1.220491e-16, 1.220584e-16, 1.220824e-16, 1.220659e-16, 1.220725e-16, 
    1.220566e-16, 1.220468e-16, 1.220516e-16, 1.220214e-16, 1.220332e-16, 
    1.21972e-16, 1.219983e-16, 1.21929e-16, 1.219455e-16, 1.21925e-16, 
    1.219354e-16, 1.219177e-16, 1.219336e-16, 1.219059e-16, 1.219e-16, 
    1.219041e-16, 1.218881e-16, 1.219345e-16, 1.219168e-16, 1.220518e-16, 
    1.22051e-16, 1.220472e-16, 1.220639e-16, 1.220648e-16, 1.220797e-16, 
    1.220663e-16, 1.220608e-16, 1.220461e-16, 1.220377e-16, 1.220296e-16, 
    1.220119e-16, 1.219923e-16, 1.219646e-16, 1.219444e-16, 1.21931e-16, 
    1.219392e-16, 1.21932e-16, 1.219401e-16, 1.219438e-16, 1.219023e-16, 
    1.219257e-16, 1.218904e-16, 1.218923e-16, 1.219084e-16, 1.218921e-16, 
    1.220505e-16, 1.22055e-16, 1.220711e-16, 1.220585e-16, 1.220813e-16, 
    1.220687e-16, 1.220616e-16, 1.220333e-16, 1.220267e-16, 1.220211e-16, 
    1.220097e-16, 1.219952e-16, 1.219699e-16, 1.219477e-16, 1.219273e-16, 
    1.219288e-16, 1.219283e-16, 1.219239e-16, 1.21935e-16, 1.21922e-16, 
    1.2192e-16, 1.219255e-16, 1.218925e-16, 1.219019e-16, 1.218923e-16, 
    1.218984e-16, 1.220535e-16, 1.220458e-16, 1.2205e-16, 1.220422e-16, 
    1.220478e-16, 1.220235e-16, 1.220162e-16, 1.219818e-16, 1.219956e-16, 
    1.219733e-16, 1.219932e-16, 1.219897e-16, 1.219732e-16, 1.21992e-16, 
    1.219492e-16, 1.219788e-16, 1.219237e-16, 1.219537e-16, 1.219218e-16, 
    1.219274e-16, 1.219181e-16, 1.219099e-16, 1.218993e-16, 1.218803e-16, 
    1.218846e-16, 1.218685e-16, 1.220343e-16, 1.220245e-16, 1.220251e-16, 
    1.220147e-16, 1.22007e-16, 1.219902e-16, 1.219635e-16, 1.219734e-16, 
    1.219549e-16, 1.219512e-16, 1.219793e-16, 1.219623e-16, 1.220178e-16, 
    1.220091e-16, 1.220141e-16, 1.220337e-16, 1.219715e-16, 1.220035e-16, 
    1.219442e-16, 1.219614e-16, 1.219111e-16, 1.219364e-16, 1.218871e-16, 
    1.218668e-16, 1.218464e-16, 1.218242e-16, 1.220189e-16, 1.220255e-16, 
    1.220134e-16, 1.21997e-16, 1.219811e-16, 1.219604e-16, 1.219582e-16, 
    1.219544e-16, 1.219442e-16, 1.219358e-16, 1.219534e-16, 1.219337e-16, 
    1.220076e-16, 1.219686e-16, 1.220283e-16, 1.220107e-16, 1.219979e-16, 
    1.220032e-16, 1.219745e-16, 1.219678e-16, 1.219408e-16, 1.219546e-16, 
    1.21872e-16, 1.219085e-16, 1.218064e-16, 1.21835e-16, 1.220279e-16, 
    1.220188e-16, 1.219873e-16, 1.220022e-16, 1.219589e-16, 1.219484e-16, 
    1.219396e-16, 1.219288e-16, 1.219275e-16, 1.21921e-16, 1.219316e-16, 
    1.219214e-16, 1.219604e-16, 1.219429e-16, 1.219906e-16, 1.219791e-16, 
    1.219843e-16, 1.219902e-16, 1.21972e-16, 1.219532e-16, 1.219524e-16, 
    1.219464e-16, 1.219304e-16, 1.219587e-16, 1.218681e-16, 1.219247e-16, 
    1.220088e-16, 1.219918e-16, 1.219888e-16, 1.219955e-16, 1.219495e-16, 
    1.219662e-16, 1.219211e-16, 1.219332e-16, 1.219133e-16, 1.219232e-16, 
    1.219247e-16, 1.219373e-16, 1.219453e-16, 1.219655e-16, 1.219818e-16, 
    1.219945e-16, 1.219915e-16, 1.219775e-16, 1.21952e-16, 1.219275e-16, 
    1.219329e-16, 1.219148e-16, 1.219621e-16, 1.219424e-16, 1.219502e-16, 
    1.2193e-16, 1.219738e-16, 1.219378e-16, 1.219831e-16, 1.219791e-16, 
    1.219665e-16, 1.219414e-16, 1.219352e-16, 1.219294e-16, 1.219329e-16, 
    1.219513e-16, 1.219541e-16, 1.219667e-16, 1.219704e-16, 1.219799e-16, 
    1.21988e-16, 1.219807e-16, 1.219732e-16, 1.219511e-16, 1.219314e-16, 
    1.219098e-16, 1.219044e-16, 1.218804e-16, 1.219005e-16, 1.218679e-16, 
    1.218965e-16, 1.218465e-16, 1.219351e-16, 1.218965e-16, 1.219658e-16, 
    1.219582e-16, 1.219449e-16, 1.219137e-16, 1.219301e-16, 1.219107e-16, 
    1.219541e-16, 1.219773e-16, 1.219827e-16, 1.219938e-16, 1.219825e-16, 
    1.219834e-16, 1.219726e-16, 1.21976e-16, 1.219503e-16, 1.219641e-16, 
    1.219249e-16, 1.219107e-16, 1.218703e-16, 1.218459e-16, 1.218204e-16, 
    1.218094e-16, 1.21806e-16, 1.218046e-16 ;

 MEG_carene_3 =
  4.842077e-17, 4.84111e-17, 4.841294e-17, 4.840524e-17, 4.840944e-17, 
    4.840446e-17, 4.841873e-17, 4.841079e-17, 4.841581e-17, 4.841979e-17, 
    4.839058e-17, 4.840488e-17, 4.837501e-17, 4.838422e-17, 4.836087e-17, 
    4.837654e-17, 4.835768e-17, 4.836113e-17, 4.83503e-17, 4.835339e-17, 
    4.833994e-17, 4.834887e-17, 4.833269e-17, 4.834197e-17, 4.834059e-17, 
    4.83492e-17, 4.840183e-17, 4.839242e-17, 4.840242e-17, 4.840107e-17, 
    4.840164e-17, 4.840942e-17, 4.841347e-17, 4.842139e-17, 4.841991e-17, 
    4.841403e-17, 4.840046e-17, 4.840494e-17, 4.83933e-17, 4.839356e-17, 
    4.838075e-17, 4.838653e-17, 4.83649e-17, 4.8371e-17, 4.835326e-17, 
    4.835774e-17, 4.83535e-17, 4.835476e-17, 4.835348e-17, 4.836005e-17, 
    4.835724e-17, 4.836296e-17, 4.838548e-17, 4.837891e-17, 4.839862e-17, 
    4.841077e-17, 4.841841e-17, 4.842398e-17, 4.842319e-17, 4.842173e-17, 
    4.841399e-17, 4.840658e-17, 4.840098e-17, 4.839728e-17, 4.83936e-17, 
    4.838295e-17, 4.837693e-17, 4.836376e-17, 4.836598e-17, 4.83621e-17, 
    4.835818e-17, 4.835181e-17, 4.835283e-17, 4.835007e-17, 4.836209e-17, 
    4.835415e-17, 4.836729e-17, 4.836371e-17, 4.839322e-17, 4.84037e-17, 
    4.84087e-17, 4.84126e-17, 4.84226e-17, 4.841573e-17, 4.841845e-17, 
    4.841185e-17, 4.840775e-17, 4.840975e-17, 4.839718e-17, 4.840208e-17, 
    4.837657e-17, 4.838754e-17, 4.835864e-17, 4.836551e-17, 4.835697e-17, 
    4.836129e-17, 4.835393e-17, 4.836055e-17, 4.834899e-17, 4.834654e-17, 
    4.834823e-17, 4.834156e-17, 4.836094e-17, 4.835356e-17, 4.840984e-17, 
    4.840951e-17, 4.840794e-17, 4.841488e-17, 4.841527e-17, 4.842146e-17, 
    4.84159e-17, 4.841358e-17, 4.840746e-17, 4.840396e-17, 4.840059e-17, 
    4.839319e-17, 4.838503e-17, 4.837347e-17, 4.836507e-17, 4.835948e-17, 
    4.836287e-17, 4.835988e-17, 4.836324e-17, 4.836479e-17, 4.83475e-17, 
    4.835725e-17, 4.834252e-17, 4.834331e-17, 4.835002e-17, 4.834322e-17, 
    4.840928e-17, 4.841115e-17, 4.841788e-17, 4.841261e-17, 4.842212e-17, 
    4.841688e-17, 4.841391e-17, 4.840212e-17, 4.839938e-17, 4.839704e-17, 
    4.839227e-17, 4.838623e-17, 4.837569e-17, 4.836644e-17, 4.835792e-17, 
    4.835854e-17, 4.835833e-17, 4.835649e-17, 4.836112e-17, 4.835572e-17, 
    4.835487e-17, 4.835718e-17, 4.834342e-17, 4.834734e-17, 4.834333e-17, 
    4.834586e-17, 4.841053e-17, 4.840734e-17, 4.840907e-17, 4.840585e-17, 
    4.840816e-17, 4.839804e-17, 4.8395e-17, 4.838066e-17, 4.838639e-17, 
    4.83771e-17, 4.838539e-17, 4.838396e-17, 4.837706e-17, 4.83849e-17, 
    4.836707e-17, 4.837939e-17, 4.835642e-17, 4.836894e-17, 4.835565e-17, 
    4.835796e-17, 4.835407e-17, 4.835066e-17, 4.834625e-17, 4.833831e-17, 
    4.834012e-17, 4.833339e-17, 4.840253e-17, 4.839846e-17, 4.83987e-17, 
    4.839436e-17, 4.839118e-17, 4.838414e-17, 4.837301e-17, 4.837715e-17, 
    4.836942e-17, 4.83679e-17, 4.837959e-17, 4.837252e-17, 4.839564e-17, 
    4.839202e-17, 4.83941e-17, 4.840228e-17, 4.837636e-17, 4.838972e-17, 
    4.836495e-17, 4.837215e-17, 4.835116e-17, 4.83617e-17, 4.834114e-17, 
    4.833268e-17, 4.83242e-17, 4.831492e-17, 4.839611e-17, 4.839889e-17, 
    4.839381e-17, 4.838701e-17, 4.838036e-17, 4.837174e-17, 4.837079e-17, 
    4.836921e-17, 4.836497e-17, 4.836147e-17, 4.836882e-17, 4.836058e-17, 
    4.839141e-17, 4.837515e-17, 4.840004e-17, 4.83927e-17, 4.838735e-17, 
    4.838958e-17, 4.83776e-17, 4.837482e-17, 4.836357e-17, 4.836932e-17, 
    4.833487e-17, 4.835009e-17, 4.830749e-17, 4.831943e-17, 4.839989e-17, 
    4.839606e-17, 4.838295e-17, 4.838917e-17, 4.83711e-17, 4.836671e-17, 
    4.836304e-17, 4.835855e-17, 4.835798e-17, 4.835531e-17, 4.83597e-17, 
    4.835544e-17, 4.837172e-17, 4.836442e-17, 4.838431e-17, 4.837953e-17, 
    4.838168e-17, 4.838414e-17, 4.837658e-17, 4.836874e-17, 4.836838e-17, 
    4.836589e-17, 4.835924e-17, 4.837102e-17, 4.833325e-17, 4.835685e-17, 
    4.839191e-17, 4.838481e-17, 4.838357e-17, 4.838636e-17, 4.836716e-17, 
    4.837413e-17, 4.835535e-17, 4.836038e-17, 4.83521e-17, 4.835622e-17, 
    4.835684e-17, 4.836211e-17, 4.836544e-17, 4.837385e-17, 4.838064e-17, 
    4.838593e-17, 4.838469e-17, 4.837887e-17, 4.836821e-17, 4.835802e-17, 
    4.836027e-17, 4.835272e-17, 4.837241e-17, 4.836424e-17, 4.836746e-17, 
    4.835904e-17, 4.83773e-17, 4.836231e-17, 4.838121e-17, 4.837951e-17, 
    4.837427e-17, 4.836381e-17, 4.836122e-17, 4.83588e-17, 4.836026e-17, 
    4.836791e-17, 4.836908e-17, 4.837435e-17, 4.83759e-17, 4.837987e-17, 
    4.838324e-17, 4.83802e-17, 4.837705e-17, 4.836783e-17, 4.835962e-17, 
    4.835064e-17, 4.834836e-17, 4.833835e-17, 4.834675e-17, 4.833315e-17, 
    4.834509e-17, 4.832425e-17, 4.836116e-17, 4.834508e-17, 4.837397e-17, 
    4.83708e-17, 4.836527e-17, 4.835224e-17, 4.835908e-17, 4.835099e-17, 
    4.836911e-17, 4.837876e-17, 4.838103e-17, 4.838564e-17, 4.838092e-17, 
    4.83813e-17, 4.837679e-17, 4.837823e-17, 4.836752e-17, 4.837326e-17, 
    4.835691e-17, 4.835101e-17, 4.833416e-17, 4.832397e-17, 4.831333e-17, 
    4.830874e-17, 4.830733e-17, 4.830675e-17 ;

 MEG_ethanol =
  3.91629e-18, 3.914856e-18, 3.915128e-18, 3.913988e-18, 3.91461e-18, 
    3.913872e-18, 3.915987e-18, 3.914811e-18, 3.915554e-18, 3.916144e-18, 
    3.911814e-18, 3.913934e-18, 3.909504e-18, 3.91087e-18, 3.907407e-18, 
    3.909732e-18, 3.906934e-18, 3.907446e-18, 3.905838e-18, 3.906296e-18, 
    3.904299e-18, 3.905625e-18, 3.903221e-18, 3.904601e-18, 3.904395e-18, 
    3.905673e-18, 3.913481e-18, 3.912087e-18, 3.91357e-18, 3.91337e-18, 
    3.913454e-18, 3.914607e-18, 3.915207e-18, 3.916381e-18, 3.916163e-18, 
    3.91529e-18, 3.913279e-18, 3.913943e-18, 3.912217e-18, 3.912255e-18, 
    3.910356e-18, 3.911212e-18, 3.908005e-18, 3.908909e-18, 3.906277e-18, 
    3.906942e-18, 3.906313e-18, 3.9065e-18, 3.90631e-18, 3.907284e-18, 
    3.906869e-18, 3.907718e-18, 3.911057e-18, 3.910083e-18, 3.913006e-18, 
    3.914808e-18, 3.91594e-18, 3.916765e-18, 3.916649e-18, 3.916432e-18, 
    3.915285e-18, 3.914186e-18, 3.913357e-18, 3.912807e-18, 3.912261e-18, 
    3.910683e-18, 3.909789e-18, 3.907836e-18, 3.908165e-18, 3.90759e-18, 
    3.907007e-18, 3.906062e-18, 3.906214e-18, 3.905803e-18, 3.907588e-18, 
    3.90641e-18, 3.908358e-18, 3.907827e-18, 3.912205e-18, 3.913759e-18, 
    3.9145e-18, 3.915079e-18, 3.91656e-18, 3.915543e-18, 3.915946e-18, 
    3.914967e-18, 3.914359e-18, 3.914656e-18, 3.912791e-18, 3.913519e-18, 
    3.909737e-18, 3.911363e-18, 3.907075e-18, 3.908095e-18, 3.906827e-18, 
    3.90747e-18, 3.906377e-18, 3.90736e-18, 3.905643e-18, 3.90528e-18, 
    3.90553e-18, 3.904539e-18, 3.907417e-18, 3.906322e-18, 3.914668e-18, 
    3.914621e-18, 3.914387e-18, 3.915417e-18, 3.915475e-18, 3.916392e-18, 
    3.915567e-18, 3.915224e-18, 3.914316e-18, 3.913797e-18, 3.913298e-18, 
    3.9122e-18, 3.91099e-18, 3.909275e-18, 3.90803e-18, 3.907201e-18, 
    3.907703e-18, 3.907261e-18, 3.907759e-18, 3.907989e-18, 3.905422e-18, 
    3.90687e-18, 3.904682e-18, 3.904799e-18, 3.905797e-18, 3.904786e-18, 
    3.914586e-18, 3.914864e-18, 3.915861e-18, 3.915081e-18, 3.91649e-18, 
    3.915713e-18, 3.915272e-18, 3.913524e-18, 3.913119e-18, 3.912771e-18, 
    3.912064e-18, 3.911169e-18, 3.909606e-18, 3.908234e-18, 3.90697e-18, 
    3.907061e-18, 3.907029e-18, 3.906757e-18, 3.907444e-18, 3.906643e-18, 
    3.906517e-18, 3.90686e-18, 3.904816e-18, 3.905398e-18, 3.904802e-18, 
    3.905178e-18, 3.914771e-18, 3.914298e-18, 3.914555e-18, 3.914078e-18, 
    3.914421e-18, 3.912919e-18, 3.91247e-18, 3.910342e-18, 3.911192e-18, 
    3.909815e-18, 3.911044e-18, 3.910832e-18, 3.909809e-18, 3.910972e-18, 
    3.908327e-18, 3.910153e-18, 3.906746e-18, 3.908604e-18, 3.906632e-18, 
    3.906975e-18, 3.906397e-18, 3.90589e-18, 3.905235e-18, 3.904056e-18, 
    3.904325e-18, 3.903324e-18, 3.913585e-18, 3.912982e-18, 3.913018e-18, 
    3.912374e-18, 3.911902e-18, 3.910858e-18, 3.909207e-18, 3.909822e-18, 
    3.908674e-18, 3.90845e-18, 3.910184e-18, 3.909135e-18, 3.912564e-18, 
    3.912028e-18, 3.912335e-18, 3.913548e-18, 3.909704e-18, 3.911685e-18, 
    3.908013e-18, 3.909081e-18, 3.905965e-18, 3.90753e-18, 3.904477e-18, 
    3.90322e-18, 3.901958e-18, 3.900578e-18, 3.912633e-18, 3.913045e-18, 
    3.912292e-18, 3.911283e-18, 3.910299e-18, 3.909019e-18, 3.908878e-18, 
    3.908644e-18, 3.908015e-18, 3.907496e-18, 3.908586e-18, 3.907364e-18, 
    3.911938e-18, 3.909524e-18, 3.913217e-18, 3.912127e-18, 3.911335e-18, 
    3.911665e-18, 3.909888e-18, 3.909476e-18, 3.907808e-18, 3.90866e-18, 
    3.903545e-18, 3.905807e-18, 3.899472e-18, 3.901249e-18, 3.913194e-18, 
    3.912627e-18, 3.910681e-18, 3.911604e-18, 3.908924e-18, 3.908273e-18, 
    3.907729e-18, 3.907063e-18, 3.906978e-18, 3.906582e-18, 3.907234e-18, 
    3.906601e-18, 3.909016e-18, 3.907933e-18, 3.910883e-18, 3.910174e-18, 
    3.910494e-18, 3.910858e-18, 3.909737e-18, 3.908574e-18, 3.908521e-18, 
    3.908153e-18, 3.907165e-18, 3.908912e-18, 3.903304e-18, 3.906811e-18, 
    3.91201e-18, 3.910958e-18, 3.910774e-18, 3.911187e-18, 3.90834e-18, 
    3.909374e-18, 3.906588e-18, 3.907334e-18, 3.906104e-18, 3.906717e-18, 
    3.906809e-18, 3.907591e-18, 3.908086e-18, 3.909332e-18, 3.910339e-18, 
    3.911124e-18, 3.910939e-18, 3.910077e-18, 3.908496e-18, 3.906984e-18, 
    3.907318e-18, 3.906197e-18, 3.909119e-18, 3.907907e-18, 3.908385e-18, 
    3.907135e-18, 3.909844e-18, 3.907621e-18, 3.910424e-18, 3.910172e-18, 
    3.909394e-18, 3.907844e-18, 3.907459e-18, 3.9071e-18, 3.907316e-18, 
    3.908451e-18, 3.908624e-18, 3.909407e-18, 3.909636e-18, 3.910224e-18, 
    3.910725e-18, 3.910275e-18, 3.909808e-18, 3.908439e-18, 3.907222e-18, 
    3.905887e-18, 3.90555e-18, 3.904063e-18, 3.905311e-18, 3.90329e-18, 
    3.905065e-18, 3.901966e-18, 3.907451e-18, 3.905062e-18, 3.909349e-18, 
    3.90888e-18, 3.908061e-18, 3.906126e-18, 3.90714e-18, 3.90594e-18, 
    3.908629e-18, 3.91006e-18, 3.910397e-18, 3.911081e-18, 3.910381e-18, 
    3.910437e-18, 3.909769e-18, 3.909982e-18, 3.908393e-18, 3.909245e-18, 
    3.906819e-18, 3.905943e-18, 3.903439e-18, 3.901925e-18, 3.900341e-18, 
    3.899658e-18, 3.899448e-18, 3.899361e-18 ;

 MEG_formaldehyde =
  7.832579e-19, 7.829713e-19, 7.830256e-19, 7.827976e-19, 7.82922e-19, 
    7.827743e-19, 7.831974e-19, 7.82962e-19, 7.831108e-19, 7.832288e-19, 
    7.823628e-19, 7.827868e-19, 7.819008e-19, 7.821741e-19, 7.814813e-19, 
    7.819464e-19, 7.813867e-19, 7.814892e-19, 7.811675e-19, 7.812593e-19, 
    7.808597e-19, 7.811251e-19, 7.806442e-19, 7.809201e-19, 7.80879e-19, 
    7.811347e-19, 7.826961e-19, 7.824173e-19, 7.82714e-19, 7.826738e-19, 
    7.826907e-19, 7.829213e-19, 7.830413e-19, 7.832761e-19, 7.832325e-19, 
    7.83058e-19, 7.826557e-19, 7.827886e-19, 7.824434e-19, 7.82451e-19, 
    7.820711e-19, 7.822424e-19, 7.81601e-19, 7.817818e-19, 7.812553e-19, 
    7.813884e-19, 7.812625e-19, 7.813e-19, 7.81262e-19, 7.814569e-19, 
    7.813737e-19, 7.815435e-19, 7.822114e-19, 7.820166e-19, 7.826011e-19, 
    7.829616e-19, 7.83188e-19, 7.83353e-19, 7.833297e-19, 7.832863e-19, 
    7.83057e-19, 7.828371e-19, 7.826713e-19, 7.825613e-19, 7.824522e-19, 
    7.821365e-19, 7.819578e-19, 7.815671e-19, 7.816329e-19, 7.815179e-19, 
    7.814014e-19, 7.812124e-19, 7.812427e-19, 7.811606e-19, 7.815175e-19, 
    7.812819e-19, 7.816716e-19, 7.815655e-19, 7.82441e-19, 7.827518e-19, 
    7.829e-19, 7.830158e-19, 7.833121e-19, 7.831085e-19, 7.831892e-19, 
    7.829935e-19, 7.828718e-19, 7.829312e-19, 7.825583e-19, 7.827038e-19, 
    7.819473e-19, 7.822726e-19, 7.81415e-19, 7.81619e-19, 7.813655e-19, 
    7.814939e-19, 7.812753e-19, 7.81472e-19, 7.811285e-19, 7.810559e-19, 
    7.811059e-19, 7.809078e-19, 7.814833e-19, 7.812643e-19, 7.829336e-19, 
    7.829241e-19, 7.828774e-19, 7.830833e-19, 7.830949e-19, 7.832783e-19, 
    7.831134e-19, 7.830447e-19, 7.828633e-19, 7.827595e-19, 7.826595e-19, 
    7.8244e-19, 7.82198e-19, 7.81855e-19, 7.81606e-19, 7.814402e-19, 
    7.815406e-19, 7.814521e-19, 7.815518e-19, 7.815977e-19, 7.810843e-19, 
    7.813739e-19, 7.809363e-19, 7.809598e-19, 7.811593e-19, 7.809571e-19, 
    7.829171e-19, 7.829728e-19, 7.831722e-19, 7.830161e-19, 7.83298e-19, 
    7.831425e-19, 7.830544e-19, 7.827049e-19, 7.826236e-19, 7.825542e-19, 
    7.824128e-19, 7.822338e-19, 7.819212e-19, 7.816467e-19, 7.813939e-19, 
    7.814121e-19, 7.814058e-19, 7.813513e-19, 7.814889e-19, 7.813285e-19, 
    7.813034e-19, 7.813719e-19, 7.809631e-19, 7.810796e-19, 7.809603e-19, 
    7.810357e-19, 7.829542e-19, 7.828597e-19, 7.82911e-19, 7.828155e-19, 
    7.828842e-19, 7.825838e-19, 7.824938e-19, 7.820684e-19, 7.822383e-19, 
    7.819629e-19, 7.822089e-19, 7.821663e-19, 7.819616e-19, 7.821943e-19, 
    7.816654e-19, 7.820307e-19, 7.813492e-19, 7.817207e-19, 7.813263e-19, 
    7.81395e-19, 7.812794e-19, 7.81178e-19, 7.81047e-19, 7.808111e-19, 
    7.808649e-19, 7.806648e-19, 7.827171e-19, 7.825963e-19, 7.826035e-19, 
    7.824748e-19, 7.823804e-19, 7.821716e-19, 7.818414e-19, 7.819643e-19, 
    7.817348e-19, 7.8169e-19, 7.820367e-19, 7.81827e-19, 7.825129e-19, 
    7.824055e-19, 7.824669e-19, 7.827095e-19, 7.819408e-19, 7.82337e-19, 
    7.816026e-19, 7.818161e-19, 7.811929e-19, 7.81506e-19, 7.808954e-19, 
    7.806439e-19, 7.803916e-19, 7.801156e-19, 7.825267e-19, 7.826091e-19, 
    7.824584e-19, 7.822566e-19, 7.820597e-19, 7.818038e-19, 7.817756e-19, 
    7.817287e-19, 7.81603e-19, 7.814991e-19, 7.817172e-19, 7.814728e-19, 
    7.823875e-19, 7.819049e-19, 7.826434e-19, 7.824254e-19, 7.82267e-19, 
    7.823329e-19, 7.819776e-19, 7.818952e-19, 7.815617e-19, 7.81732e-19, 
    7.807089e-19, 7.811613e-19, 7.798944e-19, 7.802498e-19, 7.826387e-19, 
    7.825253e-19, 7.821362e-19, 7.823207e-19, 7.817848e-19, 7.816546e-19, 
    7.815459e-19, 7.814126e-19, 7.813957e-19, 7.813163e-19, 7.814468e-19, 
    7.813202e-19, 7.818031e-19, 7.815866e-19, 7.821765e-19, 7.820348e-19, 
    7.820988e-19, 7.821715e-19, 7.819475e-19, 7.817147e-19, 7.817041e-19, 
    7.816305e-19, 7.81433e-19, 7.817825e-19, 7.806608e-19, 7.813622e-19, 
    7.824021e-19, 7.821916e-19, 7.821548e-19, 7.822375e-19, 7.816679e-19, 
    7.818748e-19, 7.813175e-19, 7.814667e-19, 7.812209e-19, 7.813434e-19, 
    7.813618e-19, 7.815181e-19, 7.816171e-19, 7.818663e-19, 7.820678e-19, 
    7.822247e-19, 7.821878e-19, 7.820153e-19, 7.816991e-19, 7.813967e-19, 
    7.814636e-19, 7.812395e-19, 7.818238e-19, 7.815814e-19, 7.816768e-19, 
    7.81427e-19, 7.819688e-19, 7.815241e-19, 7.820846e-19, 7.820343e-19, 
    7.818788e-19, 7.815687e-19, 7.814919e-19, 7.814199e-19, 7.814632e-19, 
    7.816901e-19, 7.817249e-19, 7.818813e-19, 7.819273e-19, 7.820448e-19, 
    7.821449e-19, 7.820549e-19, 7.819615e-19, 7.816877e-19, 7.814443e-19, 
    7.811774e-19, 7.8111e-19, 7.808125e-19, 7.810621e-19, 7.80658e-19, 
    7.810129e-19, 7.803931e-19, 7.814901e-19, 7.810124e-19, 7.818699e-19, 
    7.81776e-19, 7.816121e-19, 7.812251e-19, 7.814281e-19, 7.81188e-19, 
    7.817258e-19, 7.820121e-19, 7.820793e-19, 7.822162e-19, 7.820762e-19, 
    7.820873e-19, 7.819537e-19, 7.819963e-19, 7.816786e-19, 7.818489e-19, 
    7.813637e-19, 7.811885e-19, 7.806877e-19, 7.803849e-19, 7.800683e-19, 
    7.799315e-19, 7.798895e-19, 7.798722e-19 ;

 MEG_isoprene =
  6.252618e-19, 6.249929e-19, 6.250438e-19, 6.2483e-19, 6.249466e-19, 
    6.248081e-19, 6.25205e-19, 6.249842e-19, 6.251238e-19, 6.252345e-19, 
    6.24422e-19, 6.248198e-19, 6.239885e-19, 6.242449e-19, 6.235949e-19, 
    6.240313e-19, 6.235061e-19, 6.236023e-19, 6.233004e-19, 6.233865e-19, 
    6.230115e-19, 6.232605e-19, 6.228093e-19, 6.230682e-19, 6.230296e-19, 
    6.232696e-19, 6.247348e-19, 6.244731e-19, 6.247515e-19, 6.247138e-19, 
    6.247296e-19, 6.24946e-19, 6.250586e-19, 6.252789e-19, 6.25238e-19, 
    6.250742e-19, 6.246968e-19, 6.248215e-19, 6.244976e-19, 6.245047e-19, 
    6.241483e-19, 6.24309e-19, 6.237072e-19, 6.238769e-19, 6.233829e-19, 
    6.235077e-19, 6.233896e-19, 6.234247e-19, 6.233891e-19, 6.23572e-19, 
    6.234939e-19, 6.236533e-19, 6.242799e-19, 6.240972e-19, 6.246455e-19, 
    6.249838e-19, 6.251962e-19, 6.25351e-19, 6.253291e-19, 6.252884e-19, 
    6.250734e-19, 6.24867e-19, 6.247114e-19, 6.246082e-19, 6.245059e-19, 
    6.242097e-19, 6.24042e-19, 6.236754e-19, 6.237372e-19, 6.236292e-19, 
    6.235199e-19, 6.233425e-19, 6.23371e-19, 6.232939e-19, 6.236289e-19, 
    6.234077e-19, 6.237734e-19, 6.236739e-19, 6.244954e-19, 6.24787e-19, 
    6.249261e-19, 6.250347e-19, 6.253126e-19, 6.251216e-19, 6.251973e-19, 
    6.250136e-19, 6.248995e-19, 6.249552e-19, 6.246054e-19, 6.24742e-19, 
    6.240321e-19, 6.243373e-19, 6.235327e-19, 6.237241e-19, 6.234862e-19, 
    6.236067e-19, 6.234016e-19, 6.235861e-19, 6.232638e-19, 6.231957e-19, 
    6.232426e-19, 6.230566e-19, 6.235968e-19, 6.233912e-19, 6.249576e-19, 
    6.249487e-19, 6.249048e-19, 6.25098e-19, 6.251089e-19, 6.252809e-19, 
    6.251262e-19, 6.250618e-19, 6.248915e-19, 6.247941e-19, 6.247004e-19, 
    6.244944e-19, 6.242674e-19, 6.239456e-19, 6.237119e-19, 6.235564e-19, 
    6.236505e-19, 6.235675e-19, 6.23661e-19, 6.237041e-19, 6.232223e-19, 
    6.234942e-19, 6.230834e-19, 6.231055e-19, 6.232927e-19, 6.23103e-19, 
    6.24942e-19, 6.249943e-19, 6.251814e-19, 6.250349e-19, 6.252994e-19, 
    6.251535e-19, 6.250709e-19, 6.247429e-19, 6.246667e-19, 6.246016e-19, 
    6.244689e-19, 6.243009e-19, 6.240076e-19, 6.237501e-19, 6.235128e-19, 
    6.235299e-19, 6.23524e-19, 6.234729e-19, 6.23602e-19, 6.234515e-19, 
    6.234279e-19, 6.234922e-19, 6.231085e-19, 6.232178e-19, 6.23106e-19, 
    6.231767e-19, 6.249768e-19, 6.248882e-19, 6.249363e-19, 6.248467e-19, 
    6.249112e-19, 6.246294e-19, 6.245449e-19, 6.241458e-19, 6.243052e-19, 
    6.240468e-19, 6.242776e-19, 6.242376e-19, 6.240456e-19, 6.242639e-19, 
    6.237676e-19, 6.241104e-19, 6.234709e-19, 6.238196e-19, 6.234494e-19, 
    6.235139e-19, 6.234054e-19, 6.233103e-19, 6.231874e-19, 6.229658e-19, 
    6.230164e-19, 6.228286e-19, 6.247544e-19, 6.246411e-19, 6.246478e-19, 
    6.24527e-19, 6.244384e-19, 6.242426e-19, 6.239328e-19, 6.240482e-19, 
    6.238328e-19, 6.237907e-19, 6.24116e-19, 6.239193e-19, 6.245628e-19, 
    6.244621e-19, 6.245197e-19, 6.247473e-19, 6.24026e-19, 6.243978e-19, 
    6.237087e-19, 6.23909e-19, 6.233243e-19, 6.236181e-19, 6.23045e-19, 
    6.228089e-19, 6.225721e-19, 6.223129e-19, 6.245757e-19, 6.24653e-19, 
    6.245117e-19, 6.243224e-19, 6.241376e-19, 6.238975e-19, 6.23871e-19, 
    6.238271e-19, 6.237091e-19, 6.236116e-19, 6.238162e-19, 6.235869e-19, 
    6.244452e-19, 6.239923e-19, 6.246852e-19, 6.244807e-19, 6.24332e-19, 
    6.24394e-19, 6.240605e-19, 6.239832e-19, 6.236703e-19, 6.238301e-19, 
    6.2287e-19, 6.232947e-19, 6.221053e-19, 6.22439e-19, 6.246809e-19, 
    6.245745e-19, 6.242094e-19, 6.243824e-19, 6.238797e-19, 6.237575e-19, 
    6.236555e-19, 6.235304e-19, 6.235145e-19, 6.234401e-19, 6.235625e-19, 
    6.234437e-19, 6.238969e-19, 6.236937e-19, 6.242472e-19, 6.241142e-19, 
    6.241743e-19, 6.242426e-19, 6.240323e-19, 6.238139e-19, 6.23804e-19, 
    6.237349e-19, 6.235496e-19, 6.238775e-19, 6.228248e-19, 6.234831e-19, 
    6.244588e-19, 6.242614e-19, 6.242268e-19, 6.243044e-19, 6.2377e-19, 
    6.239641e-19, 6.234412e-19, 6.235812e-19, 6.233504e-19, 6.234655e-19, 
    6.234827e-19, 6.236295e-19, 6.237223e-19, 6.239562e-19, 6.241452e-19, 
    6.242925e-19, 6.242578e-19, 6.240959e-19, 6.237993e-19, 6.235155e-19, 
    6.235783e-19, 6.233679e-19, 6.239162e-19, 6.236888e-19, 6.237784e-19, 
    6.235439e-19, 6.240524e-19, 6.236351e-19, 6.24161e-19, 6.241138e-19, 
    6.239679e-19, 6.236769e-19, 6.236048e-19, 6.235373e-19, 6.235779e-19, 
    6.237908e-19, 6.238234e-19, 6.239702e-19, 6.240133e-19, 6.241236e-19, 
    6.242175e-19, 6.241331e-19, 6.240455e-19, 6.237886e-19, 6.235601e-19, 
    6.233097e-19, 6.232464e-19, 6.229672e-19, 6.232015e-19, 6.228221e-19, 
    6.231553e-19, 6.225735e-19, 6.236032e-19, 6.231548e-19, 6.239595e-19, 
    6.238714e-19, 6.237176e-19, 6.233545e-19, 6.23545e-19, 6.233197e-19, 
    6.238243e-19, 6.240929e-19, 6.24156e-19, 6.242845e-19, 6.241531e-19, 
    6.241635e-19, 6.240382e-19, 6.240781e-19, 6.2378e-19, 6.239399e-19, 
    6.234845e-19, 6.233201e-19, 6.228501e-19, 6.225658e-19, 6.222685e-19, 
    6.221402e-19, 6.221007e-19, 6.220844e-19 ;

 MEG_methanol =
  8.573229e-17, 8.571758e-17, 8.572036e-17, 8.570866e-17, 8.571505e-17, 
    8.570747e-17, 8.572918e-17, 8.57171e-17, 8.572474e-17, 8.57308e-17, 
    8.568636e-17, 8.570811e-17, 8.566265e-17, 8.567667e-17, 8.564113e-17, 
    8.566498e-17, 8.563628e-17, 8.564153e-17, 8.562505e-17, 8.562975e-17, 
    8.560928e-17, 8.562287e-17, 8.559826e-17, 8.561238e-17, 8.561028e-17, 
    8.562337e-17, 8.570346e-17, 8.568915e-17, 8.570438e-17, 8.570231e-17, 
    8.570318e-17, 8.571502e-17, 8.572117e-17, 8.573323e-17, 8.573098e-17, 
    8.572202e-17, 8.570138e-17, 8.57082e-17, 8.569049e-17, 8.569088e-17, 
    8.567139e-17, 8.568018e-17, 8.564727e-17, 8.565655e-17, 8.562955e-17, 
    8.563637e-17, 8.562992e-17, 8.563183e-17, 8.562989e-17, 8.563987e-17, 
    8.563561e-17, 8.564432e-17, 8.567859e-17, 8.566859e-17, 8.569858e-17, 
    8.571707e-17, 8.57287e-17, 8.573717e-17, 8.573597e-17, 8.573375e-17, 
    8.572198e-17, 8.571069e-17, 8.570218e-17, 8.569654e-17, 8.569094e-17, 
    8.567474e-17, 8.566557e-17, 8.564553e-17, 8.56489e-17, 8.5643e-17, 
    8.563703e-17, 8.562735e-17, 8.56289e-17, 8.562469e-17, 8.564299e-17, 
    8.563091e-17, 8.56509e-17, 8.564545e-17, 8.569036e-17, 8.570631e-17, 
    8.571392e-17, 8.571987e-17, 8.573507e-17, 8.572462e-17, 8.572876e-17, 
    8.571872e-17, 8.571247e-17, 8.571552e-17, 8.569639e-17, 8.570385e-17, 
    8.566503e-17, 8.568172e-17, 8.563773e-17, 8.564819e-17, 8.563519e-17, 
    8.564177e-17, 8.563057e-17, 8.564065e-17, 8.562305e-17, 8.561933e-17, 
    8.56219e-17, 8.561175e-17, 8.564123e-17, 8.563001e-17, 8.571564e-17, 
    8.571515e-17, 8.571276e-17, 8.572333e-17, 8.572392e-17, 8.573333e-17, 
    8.572487e-17, 8.572135e-17, 8.571203e-17, 8.57067e-17, 8.570158e-17, 
    8.569032e-17, 8.56779e-17, 8.56603e-17, 8.564752e-17, 8.563902e-17, 
    8.564417e-17, 8.563963e-17, 8.564474e-17, 8.564709e-17, 8.562079e-17, 
    8.563563e-17, 8.561321e-17, 8.561441e-17, 8.562463e-17, 8.561428e-17, 
    8.57148e-17, 8.571766e-17, 8.572789e-17, 8.571988e-17, 8.573435e-17, 
    8.572636e-17, 8.572185e-17, 8.570391e-17, 8.569974e-17, 8.569618e-17, 
    8.568892e-17, 8.567974e-17, 8.566369e-17, 8.564961e-17, 8.563665e-17, 
    8.563758e-17, 8.563726e-17, 8.563446e-17, 8.564152e-17, 8.56333e-17, 
    8.563201e-17, 8.563552e-17, 8.561458e-17, 8.562055e-17, 8.561444e-17, 
    8.56183e-17, 8.57167e-17, 8.571185e-17, 8.571449e-17, 8.570958e-17, 
    8.571311e-17, 8.569769e-17, 8.569308e-17, 8.567125e-17, 8.567997e-17, 
    8.566584e-17, 8.567845e-17, 8.567627e-17, 8.566577e-17, 8.567771e-17, 
    8.565056e-17, 8.566931e-17, 8.563436e-17, 8.565341e-17, 8.563318e-17, 
    8.563671e-17, 8.563078e-17, 8.562559e-17, 8.561888e-17, 8.560679e-17, 
    8.560955e-17, 8.559931e-17, 8.570453e-17, 8.569833e-17, 8.56987e-17, 
    8.56921e-17, 8.568726e-17, 8.567655e-17, 8.56596e-17, 8.566591e-17, 
    8.565414e-17, 8.565184e-17, 8.566962e-17, 8.565887e-17, 8.569405e-17, 
    8.568855e-17, 8.56917e-17, 8.570414e-17, 8.56647e-17, 8.568503e-17, 
    8.564735e-17, 8.56583e-17, 8.562635e-17, 8.56424e-17, 8.561112e-17, 
    8.559824e-17, 8.558533e-17, 8.557122e-17, 8.569477e-17, 8.569899e-17, 
    8.569127e-17, 8.568091e-17, 8.56708e-17, 8.565767e-17, 8.565623e-17, 
    8.565382e-17, 8.564737e-17, 8.564204e-17, 8.565324e-17, 8.564069e-17, 
    8.568762e-17, 8.566286e-17, 8.570075e-17, 8.568957e-17, 8.568144e-17, 
    8.568483e-17, 8.566659e-17, 8.566236e-17, 8.564525e-17, 8.5654e-17, 
    8.560157e-17, 8.562473e-17, 8.555992e-17, 8.557808e-17, 8.570051e-17, 
    8.569469e-17, 8.567473e-17, 8.56842e-17, 8.56567e-17, 8.565001e-17, 
    8.564444e-17, 8.563761e-17, 8.563674e-17, 8.563268e-17, 8.563936e-17, 
    8.563287e-17, 8.565764e-17, 8.564653e-17, 8.56768e-17, 8.566953e-17, 
    8.567281e-17, 8.567654e-17, 8.566504e-17, 8.56531e-17, 8.565257e-17, 
    8.564878e-17, 8.563864e-17, 8.565658e-17, 8.55991e-17, 8.563502e-17, 
    8.568837e-17, 8.567757e-17, 8.567568e-17, 8.567993e-17, 8.565071e-17, 
    8.566132e-17, 8.563273e-17, 8.564038e-17, 8.562778e-17, 8.563406e-17, 
    8.5635e-17, 8.564302e-17, 8.564809e-17, 8.566088e-17, 8.567122e-17, 
    8.567928e-17, 8.567738e-17, 8.566852e-17, 8.56523e-17, 8.563679e-17, 
    8.564022e-17, 8.562874e-17, 8.565869e-17, 8.564625e-17, 8.565116e-17, 
    8.563835e-17, 8.566614e-17, 8.564332e-17, 8.567208e-17, 8.56695e-17, 
    8.566152e-17, 8.564561e-17, 8.564167e-17, 8.563798e-17, 8.56402e-17, 
    8.565184e-17, 8.565363e-17, 8.566165e-17, 8.566401e-17, 8.567004e-17, 
    8.567517e-17, 8.567055e-17, 8.566576e-17, 8.565173e-17, 8.563923e-17, 
    8.562555e-17, 8.56221e-17, 8.560687e-17, 8.561965e-17, 8.559895e-17, 
    8.561712e-17, 8.55854e-17, 8.564158e-17, 8.56171e-17, 8.566106e-17, 
    8.565625e-17, 8.564783e-17, 8.5628e-17, 8.56384e-17, 8.56261e-17, 
    8.565367e-17, 8.566836e-17, 8.567181e-17, 8.567884e-17, 8.567165e-17, 
    8.567222e-17, 8.566537e-17, 8.566755e-17, 8.565125e-17, 8.565999e-17, 
    8.56351e-17, 8.562612e-17, 8.560048e-17, 8.558499e-17, 8.55688e-17, 
    8.556182e-17, 8.555967e-17, 8.555878e-17 ;

 MEG_pinene_a =
  7.460867e-17, 7.459253e-17, 7.459559e-17, 7.458275e-17, 7.458976e-17, 
    7.458144e-17, 7.460527e-17, 7.459201e-17, 7.46004e-17, 7.460703e-17, 
    7.455828e-17, 7.458214e-17, 7.453228e-17, 7.454766e-17, 7.450868e-17, 
    7.453484e-17, 7.450335e-17, 7.450912e-17, 7.449104e-17, 7.449619e-17, 
    7.447373e-17, 7.448865e-17, 7.446163e-17, 7.447713e-17, 7.447482e-17, 
    7.448919e-17, 7.457705e-17, 7.456135e-17, 7.457805e-17, 7.457579e-17, 
    7.457674e-17, 7.458972e-17, 7.459648e-17, 7.46097e-17, 7.460724e-17, 
    7.459742e-17, 7.457477e-17, 7.458225e-17, 7.456282e-17, 7.456325e-17, 
    7.454186e-17, 7.455151e-17, 7.451541e-17, 7.452559e-17, 7.449597e-17, 
    7.450345e-17, 7.449638e-17, 7.449848e-17, 7.449635e-17, 7.45073e-17, 
    7.450262e-17, 7.451218e-17, 7.454976e-17, 7.45388e-17, 7.45717e-17, 
    7.459198e-17, 7.460474e-17, 7.461403e-17, 7.461272e-17, 7.461028e-17, 
    7.459736e-17, 7.458498e-17, 7.457565e-17, 7.456946e-17, 7.456332e-17, 
    7.454554e-17, 7.453548e-17, 7.45135e-17, 7.451721e-17, 7.451073e-17, 
    7.450418e-17, 7.449356e-17, 7.449526e-17, 7.449064e-17, 7.451071e-17, 
    7.449746e-17, 7.451939e-17, 7.451341e-17, 7.456268e-17, 7.458018e-17, 
    7.458852e-17, 7.459504e-17, 7.461172e-17, 7.460026e-17, 7.46048e-17, 
    7.459378e-17, 7.458694e-17, 7.459028e-17, 7.456929e-17, 7.457748e-17, 
    7.45349e-17, 7.455321e-17, 7.450495e-17, 7.451642e-17, 7.450217e-17, 
    7.450939e-17, 7.44971e-17, 7.450815e-17, 7.448885e-17, 7.448476e-17, 
    7.448757e-17, 7.447644e-17, 7.450879e-17, 7.449647e-17, 7.459042e-17, 
    7.458988e-17, 7.458725e-17, 7.459884e-17, 7.45995e-17, 7.460982e-17, 
    7.460053e-17, 7.459667e-17, 7.458645e-17, 7.458061e-17, 7.457498e-17, 
    7.456263e-17, 7.454901e-17, 7.452971e-17, 7.451569e-17, 7.450637e-17, 
    7.451201e-17, 7.450704e-17, 7.451264e-17, 7.451522e-17, 7.448636e-17, 
    7.450264e-17, 7.447804e-17, 7.447936e-17, 7.449057e-17, 7.447921e-17, 
    7.458948e-17, 7.459262e-17, 7.460385e-17, 7.459505e-17, 7.461093e-17, 
    7.460218e-17, 7.459721e-17, 7.457753e-17, 7.457297e-17, 7.456906e-17, 
    7.45611e-17, 7.455102e-17, 7.453343e-17, 7.451798e-17, 7.450376e-17, 
    7.450479e-17, 7.450443e-17, 7.450137e-17, 7.45091e-17, 7.450009e-17, 
    7.449867e-17, 7.450252e-17, 7.447955e-17, 7.448609e-17, 7.447939e-17, 
    7.448362e-17, 7.459157e-17, 7.458625e-17, 7.458914e-17, 7.458376e-17, 
    7.458763e-17, 7.457072e-17, 7.456566e-17, 7.454171e-17, 7.455127e-17, 
    7.453578e-17, 7.454962e-17, 7.454722e-17, 7.45357e-17, 7.454881e-17, 
    7.451903e-17, 7.453959e-17, 7.450125e-17, 7.452214e-17, 7.449996e-17, 
    7.450382e-17, 7.449733e-17, 7.449162e-17, 7.448427e-17, 7.4471e-17, 
    7.447403e-17, 7.446279e-17, 7.457823e-17, 7.457142e-17, 7.457183e-17, 
    7.456459e-17, 7.455927e-17, 7.454752e-17, 7.452894e-17, 7.453586e-17, 
    7.452294e-17, 7.452042e-17, 7.453993e-17, 7.452813e-17, 7.456673e-17, 
    7.456069e-17, 7.456414e-17, 7.45778e-17, 7.453453e-17, 7.455683e-17, 
    7.451549e-17, 7.452752e-17, 7.449246e-17, 7.451007e-17, 7.447574e-17, 
    7.446161e-17, 7.444744e-17, 7.443195e-17, 7.456751e-17, 7.457215e-17, 
    7.456367e-17, 7.455231e-17, 7.454122e-17, 7.452682e-17, 7.452524e-17, 
    7.45226e-17, 7.451552e-17, 7.450968e-17, 7.452195e-17, 7.450819e-17, 
    7.455967e-17, 7.453251e-17, 7.457408e-17, 7.456181e-17, 7.455289e-17, 
    7.455661e-17, 7.45366e-17, 7.453196e-17, 7.45132e-17, 7.452279e-17, 
    7.446526e-17, 7.449068e-17, 7.441954e-17, 7.443949e-17, 7.457381e-17, 
    7.456743e-17, 7.454553e-17, 7.455591e-17, 7.452576e-17, 7.451842e-17, 
    7.451231e-17, 7.450481e-17, 7.450386e-17, 7.44994e-17, 7.450673e-17, 
    7.449962e-17, 7.452679e-17, 7.45146e-17, 7.45478e-17, 7.453983e-17, 
    7.454343e-17, 7.454752e-17, 7.453491e-17, 7.452181e-17, 7.452122e-17, 
    7.451707e-17, 7.450595e-17, 7.452562e-17, 7.446255e-17, 7.450197e-17, 
    7.456049e-17, 7.454865e-17, 7.454658e-17, 7.455123e-17, 7.451918e-17, 
    7.453082e-17, 7.449947e-17, 7.450786e-17, 7.449403e-17, 7.450092e-17, 
    7.450195e-17, 7.451075e-17, 7.451631e-17, 7.453034e-17, 7.454168e-17, 
    7.455051e-17, 7.454844e-17, 7.453872e-17, 7.452093e-17, 7.450392e-17, 
    7.450768e-17, 7.449508e-17, 7.452795e-17, 7.45143e-17, 7.451968e-17, 
    7.450563e-17, 7.453611e-17, 7.451108e-17, 7.454263e-17, 7.453979e-17, 
    7.453104e-17, 7.451359e-17, 7.450927e-17, 7.450522e-17, 7.450766e-17, 
    7.452042e-17, 7.452238e-17, 7.453118e-17, 7.453377e-17, 7.454039e-17, 
    7.454602e-17, 7.454095e-17, 7.45357e-17, 7.45203e-17, 7.450659e-17, 
    7.449159e-17, 7.44878e-17, 7.447108e-17, 7.448511e-17, 7.44624e-17, 
    7.448233e-17, 7.444752e-17, 7.450917e-17, 7.448231e-17, 7.453054e-17, 
    7.452526e-17, 7.451603e-17, 7.449427e-17, 7.450569e-17, 7.449219e-17, 
    7.452244e-17, 7.453854e-17, 7.454233e-17, 7.455004e-17, 7.454216e-17, 
    7.454278e-17, 7.453526e-17, 7.453766e-17, 7.451978e-17, 7.452936e-17, 
    7.450206e-17, 7.449221e-17, 7.446408e-17, 7.444706e-17, 7.442929e-17, 
    7.442162e-17, 7.441926e-17, 7.441829e-17 ;

 MEG_thujene_a =
  1.797621e-18, 1.797262e-18, 1.79733e-18, 1.797045e-18, 1.7972e-18, 
    1.797016e-18, 1.797545e-18, 1.79725e-18, 1.797437e-18, 1.797585e-18, 
    1.7965e-18, 1.797031e-18, 1.795922e-18, 1.796264e-18, 1.795397e-18, 
    1.795979e-18, 1.795279e-18, 1.795407e-18, 1.795005e-18, 1.79512e-18, 
    1.79462e-18, 1.794952e-18, 1.794351e-18, 1.794696e-18, 1.794644e-18, 
    1.794964e-18, 1.796918e-18, 1.796568e-18, 1.79694e-18, 1.79689e-18, 
    1.796911e-18, 1.7972e-18, 1.79735e-18, 1.797644e-18, 1.797589e-18, 
    1.797371e-18, 1.796867e-18, 1.797033e-18, 1.796601e-18, 1.796611e-18, 
    1.796135e-18, 1.79635e-18, 1.795547e-18, 1.795773e-18, 1.795115e-18, 
    1.795281e-18, 1.795124e-18, 1.795171e-18, 1.795123e-18, 1.795367e-18, 
    1.795263e-18, 1.795475e-18, 1.796311e-18, 1.796067e-18, 1.796799e-18, 
    1.79725e-18, 1.797534e-18, 1.79774e-18, 1.797711e-18, 1.797657e-18, 
    1.79737e-18, 1.797094e-18, 1.796887e-18, 1.796749e-18, 1.796612e-18, 
    1.796217e-18, 1.795993e-18, 1.795505e-18, 1.795587e-18, 1.795443e-18, 
    1.795297e-18, 1.795061e-18, 1.795099e-18, 1.794996e-18, 1.795442e-18, 
    1.795148e-18, 1.795635e-18, 1.795502e-18, 1.796598e-18, 1.796987e-18, 
    1.797173e-18, 1.797318e-18, 1.797689e-18, 1.797434e-18, 1.797535e-18, 
    1.79729e-18, 1.797138e-18, 1.797212e-18, 1.796745e-18, 1.796927e-18, 
    1.79598e-18, 1.796388e-18, 1.795314e-18, 1.795569e-18, 1.795252e-18, 
    1.795413e-18, 1.79514e-18, 1.795386e-18, 1.794956e-18, 1.794866e-18, 
    1.794928e-18, 1.79468e-18, 1.7954e-18, 1.795126e-18, 1.797215e-18, 
    1.797203e-18, 1.797145e-18, 1.797402e-18, 1.797417e-18, 1.797647e-18, 
    1.79744e-18, 1.797354e-18, 1.797127e-18, 1.796997e-18, 1.796872e-18, 
    1.796597e-18, 1.796294e-18, 1.795865e-18, 1.795553e-18, 1.795346e-18, 
    1.795471e-18, 1.795361e-18, 1.795485e-18, 1.795543e-18, 1.794901e-18, 
    1.795263e-18, 1.794716e-18, 1.794745e-18, 1.794995e-18, 1.794742e-18, 
    1.797194e-18, 1.797264e-18, 1.797514e-18, 1.797318e-18, 1.797671e-18, 
    1.797477e-18, 1.797366e-18, 1.796928e-18, 1.796827e-18, 1.79674e-18, 
    1.796563e-18, 1.796339e-18, 1.795948e-18, 1.795604e-18, 1.795288e-18, 
    1.795311e-18, 1.795303e-18, 1.795235e-18, 1.795407e-18, 1.795206e-18, 
    1.795175e-18, 1.79526e-18, 1.794749e-18, 1.794895e-18, 1.794746e-18, 
    1.79484e-18, 1.797241e-18, 1.797122e-18, 1.797187e-18, 1.797067e-18, 
    1.797153e-18, 1.796777e-18, 1.796664e-18, 1.796132e-18, 1.796345e-18, 
    1.796e-18, 1.796308e-18, 1.796255e-18, 1.795998e-18, 1.796289e-18, 
    1.795627e-18, 1.796085e-18, 1.795232e-18, 1.795697e-18, 1.795203e-18, 
    1.795289e-18, 1.795145e-18, 1.795018e-18, 1.794854e-18, 1.79456e-18, 
    1.794627e-18, 1.794377e-18, 1.796944e-18, 1.796793e-18, 1.796802e-18, 
    1.796641e-18, 1.796523e-18, 1.796261e-18, 1.795848e-18, 1.796002e-18, 
    1.795715e-18, 1.795658e-18, 1.796092e-18, 1.79583e-18, 1.796688e-18, 
    1.796554e-18, 1.796631e-18, 1.796934e-18, 1.795972e-18, 1.796468e-18, 
    1.795549e-18, 1.795816e-18, 1.795037e-18, 1.795428e-18, 1.794665e-18, 
    1.794351e-18, 1.794036e-18, 1.793691e-18, 1.796706e-18, 1.796809e-18, 
    1.79662e-18, 1.796367e-18, 1.796121e-18, 1.795801e-18, 1.795765e-18, 
    1.795707e-18, 1.795549e-18, 1.79542e-18, 1.795692e-18, 1.795387e-18, 
    1.796531e-18, 1.795927e-18, 1.796852e-18, 1.796579e-18, 1.79638e-18, 
    1.796463e-18, 1.796018e-18, 1.795915e-18, 1.795498e-18, 1.795711e-18, 
    1.794432e-18, 1.794997e-18, 1.793416e-18, 1.793859e-18, 1.796846e-18, 
    1.796704e-18, 1.796217e-18, 1.796448e-18, 1.795777e-18, 1.795614e-18, 
    1.795478e-18, 1.795311e-18, 1.79529e-18, 1.795191e-18, 1.795354e-18, 
    1.795196e-18, 1.7958e-18, 1.795529e-18, 1.796267e-18, 1.79609e-18, 
    1.79617e-18, 1.796261e-18, 1.795981e-18, 1.795689e-18, 1.795676e-18, 
    1.795584e-18, 1.795337e-18, 1.795774e-18, 1.794372e-18, 1.795248e-18, 
    1.79655e-18, 1.796286e-18, 1.79624e-18, 1.796344e-18, 1.795631e-18, 
    1.79589e-18, 1.795192e-18, 1.795379e-18, 1.795072e-18, 1.795225e-18, 
    1.795248e-18, 1.795443e-18, 1.795567e-18, 1.795879e-18, 1.796131e-18, 
    1.796328e-18, 1.796281e-18, 1.796065e-18, 1.79567e-18, 1.795291e-18, 
    1.795375e-18, 1.795095e-18, 1.795826e-18, 1.795522e-18, 1.795642e-18, 
    1.795329e-18, 1.796007e-18, 1.795451e-18, 1.796152e-18, 1.796089e-18, 
    1.795895e-18, 1.795506e-18, 1.79541e-18, 1.79532e-18, 1.795375e-18, 
    1.795659e-18, 1.795702e-18, 1.795898e-18, 1.795955e-18, 1.796103e-18, 
    1.796228e-18, 1.796115e-18, 1.795998e-18, 1.795656e-18, 1.795351e-18, 
    1.795017e-18, 1.794933e-18, 1.794561e-18, 1.794873e-18, 1.794368e-18, 
    1.794812e-18, 1.794037e-18, 1.795408e-18, 1.794811e-18, 1.795884e-18, 
    1.795766e-18, 1.795561e-18, 1.795077e-18, 1.795331e-18, 1.795031e-18, 
    1.795703e-18, 1.796061e-18, 1.796146e-18, 1.796317e-18, 1.796142e-18, 
    1.796156e-18, 1.795988e-18, 1.796042e-18, 1.795644e-18, 1.795857e-18, 
    1.79525e-18, 1.795031e-18, 1.794406e-18, 1.794027e-18, 1.793633e-18, 
    1.793462e-18, 1.793409e-18, 1.793388e-18 ;

 MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 M_LITR1C_TO_LEACHING =
  -4.065596e-25, 1.318573e-25, 2.197628e-26, 7.691677e-26, -5.521519e-25, 
    -1.565803e-25, -2.884375e-25, 3.708484e-25, -5.219339e-26, -4.120536e-25, 
    5.76876e-26, -6.318148e-26, -4.093066e-25, 2.17015e-25, -8.515768e-26, 
    2.637145e-25, 9.889298e-26, -1.922916e-25, -1.428452e-25, -3.296429e-25, 
    -4.120529e-26, -1.950387e-25, -7.416958e-26, -4.395231e-26, 
    -3.571124e-26, 1.758097e-25, -3.323899e-25, -3.900774e-25, -7.032382e-25, 
    6.043463e-26, -1.016398e-25, 9.06519e-26, -1.813036e-25, -2.389911e-25, 
    -2.197612e-26, -5.246816e-25, -2.28003e-25, 6.208277e-25, -1.813036e-25, 
    1.977859e-25, -1.593274e-25, -1.483393e-25, 1.867978e-25, 1.785567e-25, 
    -2.032798e-25, -4.56006e-25, 1.730626e-25, 2.225091e-25, -5.081995e-25, 
    -2.170149e-25, -2.142679e-25, 1.538335e-25, -1.648214e-25, -2.747016e-26, 
    -6.428037e-25, 1.428454e-25, -6.043446e-26, 1.291103e-25, -2.25256e-25, 
    -2.3075e-25, -4.58753e-25, -1.895446e-25, -4.120536e-25, -2.197612e-26, 
    -9.889281e-26, -6.043446e-26, -1.785565e-25, 5.933575e-25, -4.120529e-26, 
    2.032799e-25, 1.263632e-25, 3.18655e-25, -2.444851e-25, -4.230417e-25, 
    7.197206e-25, 1.04387e-25, 9.06519e-26, 2.362442e-25, -2.829435e-25, 
    -2.087738e-25, 3.24149e-25, -8.790471e-26, -1.867976e-25, -1.098809e-25, 
    1.428454e-25, -2.472321e-25, -2.911845e-25, -3.681012e-25, -9.339876e-26, 
    -3.571124e-26, -2.637143e-25, -6.592851e-26, 1.098811e-25, -3.818364e-25, 
    1.208692e-25, -1.23616e-25, 1.648216e-25, -7.82902e-25, -4.120529e-26, 
    -1.291101e-25, -1.730625e-25, -4.752352e-25, -5.027055e-25, 2.197628e-26, 
    -4.340298e-25, 7.691677e-26, -4.120536e-25, 1.04387e-25, 4.862235e-25, 
    2.747033e-26, -8.515768e-26, 2.939317e-25, 2.719555e-25, 1.153751e-25, 
    -2.719554e-25, -1.813036e-25, -3.296429e-25, -2.966786e-25, 
    -1.016398e-25, -1.263631e-25, -3.653542e-25, -2.966786e-25, 
    -9.614578e-26, -2.197612e-26, -7.142256e-26, -7.966364e-26, 4.010657e-25, 
    -3.104137e-25, -3.845826e-26, -1.318571e-25, 3.763425e-25, 2.197621e-25, 
    3.57114e-26, -4.669934e-26, -2.746942e-27, -5.109465e-25, -3.873304e-25, 
    1.236162e-25, -1.263631e-25, 2.444853e-25, -1.703155e-25, -3.488721e-25, 
    -1.922916e-25, 4.944653e-26, 9.339892e-26, -2.197612e-26, 4.120538e-25, 
    -3.021727e-25, 8.241083e-26, 1.785567e-25, -1.620744e-25, -9.065174e-26, 
    8.515785e-26, 2.389912e-25, 6.86757e-26, 2.060269e-25, -1.126279e-25, 
    1.703156e-25, -6.043446e-26, 4.395241e-25, 9.889298e-26, -9.614578e-26, 
    4.120545e-26, -1.813036e-25, -4.175477e-25, 9.339892e-26, -4.120529e-26, 
    3.296431e-25, -1.895446e-25, -2.582203e-25, -1.291101e-25, -5.493967e-27, 
    -1.18122e-25, -1.071339e-25, 7.416968e-25, 2.197628e-26, -1.263631e-25, 
    -7.416958e-26, -2.36244e-25, 1.867978e-25, -3.845826e-26, -7.142256e-26, 
    3.708484e-25, -7.416958e-26, 1.208692e-25, 6.86757e-26, 3.18655e-25, 
    -4.917174e-25, -1.620744e-25, -2.28003e-25, 2.389912e-25, 1.428454e-25, 
    -1.977857e-25, 1.922926e-26, -2.994256e-25, -1.922916e-25, 2.389912e-25, 
    7.691677e-26, 3.104139e-25, -3.571131e-25, 4.889705e-25, 1.455924e-25, 
    9.614595e-26, -1.098802e-26, -5.356697e-25, 3.076668e-25, -9.065174e-26, 
    -4.285358e-25, 8.241083e-26, -5.219339e-26, -2.032798e-25, 2.829436e-25, 
    -2.36244e-25, -1.922916e-25, 4.807294e-25, -1.950387e-25, 2.637145e-25, 
    8.241083e-26, 6.86757e-26, 8.241083e-26, -1.318571e-25, 3.296438e-26, 
    -8.790471e-26, -1.428452e-25, -3.681012e-25, 4.395248e-26, -1.18122e-25, 
    8.257456e-32, -4.257888e-25, 8.257438e-32, -2.170149e-25, 1.291103e-25, 
    -1.922909e-26, -5.768744e-26, -2.884375e-25, -4.395239e-25, 2.747107e-27, 
    -4.093066e-25, 1.867978e-25, -2.966786e-25, 1.318573e-25, 1.922918e-25, 
    -3.37884e-25, 1.730626e-25, 1.922926e-26, 8.515785e-26, -1.867976e-25, 
    -2.582203e-25, -5.494049e-25, -6.867554e-26, 2.911847e-25, -6.318148e-26, 
    -2.499792e-25, -1.15375e-25, 2.225091e-25, -2.3075e-25, -5.027055e-25, 
    -3.351369e-25, -3.845826e-26, -1.813036e-25, 3.543663e-25, 2.472331e-26, 
    -1.867976e-25, -2.032798e-25, 7.416975e-26, -4.53259e-25, -2.856905e-25, 
    -3.37884e-25, 1.648216e-25, -7.966364e-26, 1.483394e-25, -7.142256e-26, 
    4.395248e-26, -2.389911e-25, -5.768744e-26, -5.768744e-26, -6.867554e-26, 
    1.867978e-25, -5.494041e-26, -3.021719e-26, 1.538335e-25, 2.005329e-25, 
    5.494132e-27, -6.867554e-26, -7.966364e-26, -2.3075e-25, -5.60393e-25, 
    -9.889281e-26, -2.005327e-25, 1.236162e-25, -3.873304e-25, -2.36244e-25, 
    -9.339876e-26, 9.06519e-26, 2.747033e-26, 1.510864e-25, -4.642471e-25, 
    -2.197619e-25, -2.472321e-25, 8.790487e-26, -5.494041e-26, -5.081995e-25, 
    -1.071339e-25, 9.889298e-26, 8.241083e-26, 1.071341e-25, -2.527262e-25, 
    -3.268959e-25, -1.895446e-25, -4.53259e-25, -1.428452e-25, -3.214018e-25, 
    8.257409e-32, -2.197619e-25, -3.955715e-25, -1.263631e-25, 2.060269e-25, 
    1.236162e-25, -5.109465e-25, -1.922909e-26, 2.719555e-25, 9.889298e-26, 
    -9.889281e-26, -3.021719e-26, 3.488722e-25, -2.829435e-25, -3.955715e-25, 
    -5.081995e-25, 5.796223e-25, 9.614595e-26, -2.417381e-25, -1.977857e-25, 
    5.851164e-25, -7.142256e-26, -9.614578e-26, -3.46125e-25, 2.911847e-25, 
    1.648216e-25 ;

 M_LITR2C_TO_LEACHING =
  9.614592e-26, 6.318163e-26, 1.318572e-25, -1.016399e-25, -3.296424e-26, 
    9.889295e-26, 2.637144e-25, -4.395234e-26, 4.94465e-26, 6.867567e-26, 
    -1.455923e-25, -1.318571e-25, -1.15375e-25, 5.351441e-32, -1.043869e-25, 
    -4.862233e-25, -3.40631e-25, -3.40631e-25, 2.17015e-25, -1.922917e-25, 
    1.153751e-25, -2.362441e-25, 1.400983e-25, 4.395245e-26, 6.04346e-26, 
    4.94465e-26, -2.3075e-25, 8.790485e-26, -1.016399e-25, 3.84584e-26, 
    -5.768747e-26, -1.648214e-25, -2.499792e-25, 1.648215e-25, -3.653542e-25, 
    -3.323899e-25, 4.395245e-26, -1.263631e-25, 5.494103e-27, -3.241489e-25, 
    6.318163e-26, -3.241489e-25, 1.428453e-25, 5.768757e-26, -8.241021e-27, 
    3.955716e-25, -9.339879e-26, 4.395245e-26, 2.472328e-26, -1.043869e-25, 
    2.472323e-25, 2.307501e-25, 1.483394e-25, 2.225091e-25, -1.016399e-25, 
    4.94465e-26, 1.263632e-25, -7.691664e-26, 3.021733e-26, -3.241489e-25, 
    1.236162e-25, 1.373513e-25, -5.493996e-27, 1.126281e-25, 1.510864e-25, 
    -5.493996e-27, 9.889295e-26, -1.071339e-25, -8.515771e-26, -9.889284e-26, 
    1.922923e-26, -2.197614e-26, 2.527263e-25, -8.241069e-26, -1.538333e-25, 
    -1.098809e-25, 1.455924e-25, 2.747078e-27, 1.153751e-25, -1.098805e-26, 
    -1.648209e-26, 9.889295e-26, -6.867557e-26, -9.614581e-26, -1.648209e-26, 
    -6.318152e-26, 8.241128e-27, -1.648209e-26, 1.208691e-25, 3.296435e-26, 
    1.620745e-25, -1.428452e-25, 1.098815e-26, 2.14268e-25, -8.241069e-26, 
    -2.032798e-25, 1.181221e-25, 1.373518e-26, 1.703156e-25, 2.747078e-27, 
    -4.120537e-25, 4.94465e-26, -1.15375e-25, -2.472317e-26, -1.373512e-25, 
    1.098815e-26, 3.571138e-26, 3.296435e-26, 3.516192e-25, -8.241069e-26, 
    1.0164e-25, -9.339879e-26, -1.18122e-25, -8.241021e-27, -1.593274e-25, 
    5.494055e-26, -2.25256e-25, 2.11521e-25, 9.889295e-26, -4.944639e-26, 
    5.494055e-26, -3.845829e-26, -2.005328e-25, -3.296424e-26, 3.84584e-26, 
    -7.142259e-26, 1.0164e-25, 8.24108e-26, -1.263631e-25, 2.74703e-26, 
    -4.120532e-26, -2.746971e-27, 2.472323e-25, 5.219352e-26, 7.14227e-26, 
    -6.318152e-26, -5.494044e-26, -1.703155e-25, -3.323899e-25, 8.241128e-27, 
    3.296435e-26, 2.280031e-25, 2.19762e-25, -2.444852e-25, 2.14268e-25, 
    -5.356698e-25, -3.021727e-25, 4.395245e-26, 4.94465e-26, -3.296424e-26, 
    -2.142679e-25, 7.691675e-26, -9.065177e-26, -4.45018e-25, -1.593274e-25, 
    -4.175477e-25, -1.12628e-25, 1.703156e-25, -6.867557e-26, 6.04346e-26, 
    1.565805e-25, -1.538333e-25, 2.966787e-25, -1.977857e-25, 4.120543e-26, 
    1.09881e-25, -1.236161e-25, 3.296435e-26, 4.120543e-26, -2.664613e-25, 
    -1.813036e-25, -9.614581e-26, -1.922917e-25, 9.889295e-26, -3.049197e-25, 
    -5.493996e-27, 1.977858e-25, -2.801965e-25, 3.571138e-26, -1.098809e-25, 
    6.592865e-26, -3.186548e-25, -1.703155e-25, 1.620745e-25, -2.746971e-27, 
    -2.142679e-25, -3.845829e-26, 8.515782e-26, -1.18122e-25, 1.236162e-25, 
    -2.060268e-25, 7.14227e-26, 2.252561e-25, -7.691664e-26, 5.768757e-26, 
    2.856906e-25, 9.339889e-26, -7.142259e-26, 9.065187e-26, -1.867976e-25, 
    2.472323e-25, -1.098805e-26, 2.197625e-26, 1.922918e-25, -1.510863e-25, 
    -9.889284e-26, -2.527262e-25, 1.867977e-25, 1.09881e-25, 3.900776e-25, 
    5.351446e-32, 1.758096e-25, -1.071339e-25, 9.889295e-26, -1.922912e-26, 
    -4.669937e-26, 2.389912e-25, 3.296435e-26, -1.538333e-25, -3.296424e-26, 
    -7.966367e-26, -6.043449e-26, 1.04387e-25, 5.494103e-27, 1.098815e-26, 
    -1.236161e-25, 1.922923e-26, -2.472317e-26, 2.747078e-27, -9.339879e-26, 
    -9.339879e-26, 6.592865e-26, 5.351397e-32, -1.098805e-26, -2.74702e-26, 
    -7.966367e-26, -4.120532e-26, -6.318152e-26, -9.614581e-26, 
    -1.016399e-25, -2.746971e-27, 1.483394e-25, 5.351426e-32, -4.944639e-26, 
    -4.944639e-26, -4.944639e-26, 3.296435e-26, 1.483394e-25, -1.730625e-25, 
    -3.104137e-25, 3.29643e-25, -1.593274e-25, 3.296435e-26, -1.730625e-25, 
    5.351432e-32, -1.263631e-25, 1.840507e-25, -2.142679e-25, -4.395234e-26, 
    2.087739e-25, -2.637143e-25, 2.472323e-25, -1.538333e-25, 1.098815e-26, 
    -1.428452e-25, -1.291101e-25, -2.692084e-25, 1.318572e-25, 5.494103e-27, 
    2.362442e-25, 1.291102e-25, -1.071339e-25, -1.18122e-25, 8.24108e-26, 
    -2.142679e-25, 2.252561e-25, -1.373507e-26, -3.296424e-26, 2.060269e-25, 
    1.922918e-25, -7.142259e-26, -5.493996e-27, -1.538333e-25, -1.318571e-25, 
    -8.790474e-26, -1.922917e-25, -6.592854e-26, 1.922923e-26, -5.494044e-26, 
    3.571138e-26, 1.263632e-25, 4.395245e-26, -8.790474e-26, 9.065187e-26, 
    -1.098805e-26, -2.115208e-25, -9.339879e-26, -7.966367e-26, 
    -1.840506e-25, 1.126281e-25, 2.74703e-26, 2.197625e-26, 1.153751e-25, 
    -2.719554e-25, -2.225089e-25, -2.032798e-25, -4.944639e-26, 
    -1.373507e-26, -2.692084e-25, -1.15375e-25, -7.691664e-26, 3.461252e-25, 
    -1.538333e-25, -6.592854e-26, -1.428452e-25, -1.565804e-25, 1.04387e-25, 
    -6.043449e-26, -1.565804e-25, -1.867976e-25, -3.021722e-26, 5.351437e-32, 
    -7.691664e-26, 3.845835e-25, -7.691664e-26, -2.362441e-25, -1.346042e-25, 
    -8.241069e-26, 1.373518e-26, -1.977857e-25, -3.021727e-25, -1.20869e-25, 
    -2.25256e-25, 1.64822e-26, -6.098394e-25, 5.219352e-26, 2.334972e-25, 
    1.483394e-25 ;

 M_LITR3C_TO_LEACHING =
  2.67573e-32, -2.747022e-26, -3.021725e-26, 3.433784e-26, -6.592857e-26, 
    7.416969e-26, -4.669939e-26, -7.416964e-26, -2.472322e-25, -1.840506e-25, 
    -2.595938e-25, -5.219344e-26, -1.37351e-26, -1.098807e-26, -1.785563e-26, 
    -8.241047e-27, -7.416964e-26, 4.257891e-26, 1.813037e-25, -1.648212e-26, 
    -3.296427e-26, 1.648217e-26, -5.219344e-26, 6.592862e-26, -4.807291e-26, 
    -5.219344e-26, 3.296432e-26, 1.222426e-25, -9.61456e-27, 4.944647e-26, 
    -8.515774e-26, 1.112545e-25, -2.746998e-27, -9.20253e-26, -9.889287e-26, 
    -9.889287e-26, 8.241077e-26, -3.296427e-26, 3.02173e-26, 9.614614e-27, 
    2.747052e-27, 6.867565e-26, 2.675714e-32, -5.219344e-26, -1.208691e-25, 
    -5.768749e-26, 5.768755e-26, -1.291101e-25, 3.845837e-26, 6.592862e-26, 
    -7.00491e-26, -9.889287e-26, 1.030135e-25, -1.208691e-25, 1.263632e-25, 
    9.614589e-26, -1.648212e-26, 1.09881e-25, -6.043452e-26, -3.845832e-26, 
    -1.236161e-25, 9.614614e-27, 1.098813e-26, -4.807291e-26, 6.043457e-26, 
    -4.532588e-26, -1.057604e-25, 2.747052e-27, -3.296427e-26, 1.098813e-26, 
    -3.021725e-26, 8.241101e-27, -3.845832e-26, -3.296427e-26, -1.318572e-25, 
    1.648215e-25, 2.472325e-26, -1.922915e-26, 6.31816e-26, -2.47232e-26, 
    -2.060266e-26, -2.128944e-25, -8.790477e-26, -3.433778e-26, 2.675729e-32, 
    -6.455506e-26, 5.356701e-26, 4.257891e-26, 1.098813e-26, -4.395237e-26, 
    -7.966369e-26, 7.691672e-26, 1.455923e-25, 6.043457e-26, -1.428453e-25, 
    1.373515e-26, -3.433778e-26, 3.708486e-26, 9.202536e-26, -6.867559e-26, 
    4.120564e-27, 7.416969e-26, -1.098807e-26, 1.098813e-26, -6.730208e-26, 
    -3.021725e-26, -5.219344e-26, -1.648212e-26, 3.296432e-26, 3.159081e-26, 
    -8.241047e-27, 7.966375e-26, 1.098813e-26, 1.785566e-25, -4.532588e-26, 
    -1.483393e-25, 1.620745e-25, -4.395237e-26, -9.477233e-26, -1.208691e-25, 
    8.241101e-27, -4.395237e-26, -1.867977e-25, 6.31816e-26, 4.395242e-26, 
    8.653131e-26, 5.494076e-27, 2.334974e-26, -5.081993e-26, -3.296427e-26, 
    -1.373486e-27, 8.241077e-26, 7.142267e-26, -2.47232e-26, 9.477238e-26, 
    1.236161e-25, -4.120535e-26, 7.004916e-26, -4.120535e-26, -7.829018e-26, 
    -3.433778e-26, -5.768749e-26, 5.081998e-26, -1.799301e-25, 3.296432e-26, 
    -2.746998e-27, 5.494076e-27, -1.37351e-26, -2.334968e-26, 3.02173e-26, 
    -1.607009e-25, -3.57113e-26, -4.669939e-26, -5.219344e-26, -1.291101e-25, 
    -2.747022e-26, -5.631398e-26, 1.236164e-26, -5.631398e-26, 1.373539e-27, 
    -1.098807e-26, -1.15375e-25, -6.867559e-26, -8.241071e-26, 8.653131e-26, 
    -2.746998e-27, -9.889287e-26, -4.257886e-26, 9.202536e-26, 7.142267e-26, 
    -4.120511e-27, -1.098807e-26, -1.140015e-25, -2.884373e-26, 2.115209e-25, 
    1.222426e-25, -1.483393e-25, 1.92292e-26, -3.845832e-26, -1.648212e-26, 
    -1.318572e-25, 2.197622e-26, 5.768755e-26, -1.442188e-25, -1.15375e-25, 
    2.060271e-26, 3.296432e-26, 5.494052e-26, -2.746998e-27, -6.318154e-26, 
    4.257891e-26, 1.236164e-26, -3.845832e-26, -1.071339e-25, 1.648217e-26, 
    -1.12628e-25, 5.906106e-26, -1.043869e-25, -4.944642e-26, -8.241047e-27, 
    3.02173e-26, -1.263631e-25, -1.140015e-25, 4.12054e-26, -3.159076e-26, 
    5.768755e-26, -2.060266e-26, -1.648215e-25, -1.057604e-25, -5.631398e-26, 
    9.889292e-26, 1.373539e-27, 1.236164e-26, 2.197622e-26, 1.153751e-25, 
    1.098813e-26, 2.060271e-26, 1.675685e-25, -3.983183e-26, 7.142267e-26, 
    -3.296427e-26, 3.159081e-26, 3.708486e-26, -6.867535e-27, -4.120511e-27, 
    9.614589e-26, -2.746998e-27, 8.241101e-27, 2.747052e-27, -1.236158e-26, 
    2.609676e-26, 4.120564e-27, 1.785569e-26, -7.00491e-26, -4.944642e-26, 
    3.983189e-26, 2.747052e-27, -1.208691e-25, 6.867565e-26, 3.159081e-26, 
    -5.768749e-26, 1.098813e-26, -1.620744e-25, -6.318154e-26, -2.47232e-26, 
    -1.208691e-25, -6.180803e-26, 1.483394e-25, 1.565804e-25, -1.455923e-25, 
    -1.09881e-25, -3.57113e-26, 2.334974e-26, -1.373486e-27, 7.966375e-26, 
    -3.021725e-26, -2.197617e-26, -8.790477e-26, 5.21935e-26, 5.631404e-26, 
    -1.236161e-25, -2.747022e-26, -1.043869e-25, 9.614614e-27, 1.263632e-25, 
    -5.356696e-26, 1.648217e-26, -8.790477e-26, -9.339881e-26, -4.669939e-26, 
    1.373539e-27, 2.609676e-26, -7.691667e-26, -3.296427e-26, 6.31816e-26, 
    3.983189e-26, -7.416964e-26, -1.37351e-26, -8.241047e-27, -3.708481e-26, 
    -4.120535e-26, -6.730208e-26, 7.004916e-26, 7.829024e-26, 5.081998e-26, 
    1.497129e-25, 4.944647e-26, -4.944642e-26, -1.277366e-25, -1.922915e-26, 
    1.098813e-26, -6.730208e-26, -9.889287e-26, -3.021725e-26, -1.37351e-26, 
    -4.120535e-26, 5.768755e-26, 5.494076e-27, 8.241077e-26, 1.194956e-25, 
    7.142267e-26, -1.400982e-25, 3.159081e-26, 5.21935e-26, 2.747052e-27, 
    -6.867559e-26, 3.571135e-26, -1.922915e-26, 9.889292e-26, 2.472325e-26, 
    2.884379e-26, 3.571135e-26, 8.790482e-26, -5.219344e-26, -3.57113e-26, 
    -6.043452e-26, 1.07134e-25, -1.455923e-25, 8.515779e-26, 2.334974e-26, 
    7.142267e-26, 9.614589e-26, 1.936653e-25, -6.867559e-26, -5.219344e-26, 
    -2.747022e-26, -1.373486e-27, -1.15375e-25, 1.648217e-26, 1.703156e-25, 
    -2.747022e-26, -1.648212e-26, -2.060266e-26, -1.785563e-26, 8.241101e-27, 
    3.708486e-26, 2.005328e-25, 7.691672e-26 ;

 M_SOIL1C_TO_LEACHING =
  4.77292e-20, -1.126484e-20, -1.966279e-20, 8.172053e-21, 2.407995e-21, 
    -2.84789e-20, 2.611019e-20, 6.473118e-21, -1.506417e-20, -1.99933e-20, 
    -1.073585e-20, 7.3377e-21, 1.202228e-20, 9.449415e-21, -1.614928e-20, 
    8.778837e-22, 1.306612e-20, 7.075879e-21, -3.120186e-20, 1.089022e-20, 
    -1.361546e-20, 1.017462e-20, -2.451503e-22, -1.458524e-20, -7.966492e-21, 
    -5.315598e-21, -9.630646e-21, 7.396517e-21, 2.195094e-20, -1.979538e-20, 
    -7.422259e-21, -3.322342e-20, -9.060965e-21, 1.405001e-20, 4.959677e-21, 
    6.940484e-21, 1.540488e-20, 1.902495e-21, -1.987484e-20, 2.942888e-20, 
    -1.02586e-20, 1.615042e-20, 7.687738e-21, 4.204998e-20, 2.336374e-20, 
    9.312859e-21, -4.791148e-21, 1.449616e-20, 8.721111e-21, 2.33759e-20, 
    -1.501979e-20, -1.094535e-20, 1.012966e-20, -7.228015e-21, 8.353006e-21, 
    2.590068e-20, -4.058329e-21, -5.406638e-21, -1.333157e-20, 8.014269e-21, 
    -1.763195e-20, 2.805426e-20, 5.880907e-22, 1.204237e-20, -1.356061e-20, 
    2.083246e-20, -1.631441e-20, 2.259075e-20, 3.305067e-20, -3.941861e-20, 
    2.142675e-20, -2.516296e-21, -1.548855e-20, 2.460097e-20, -1.468248e-20, 
    -4.530471e-21, 3.332973e-20, 2.149461e-20, 4.817724e-21, -2.304878e-20, 
    3.948365e-20, -1.146841e-20, -2.936755e-20, 1.945048e-20, -3.521469e-20, 
    -1.081616e-20, 2.663862e-20, -2.051381e-20, 2.724194e-20, -5.198657e-20, 
    -3.613864e-20, 7.5427e-21, 1.245448e-21, -1.530168e-20, -2.627361e-20, 
    1.32629e-20, -2.359332e-20, 9.457282e-22, -4.267816e-21, 1.213339e-20, 
    6.413746e-21, -5.114005e-20, -5.165784e-21, 3.657119e-21, -1.052494e-20, 
    -5.089918e-20, 1.035361e-20, 1.206666e-20, 2.426423e-20, -7.814971e-21, 
    1.430281e-20, 6.451623e-21, -3.043318e-21, -8.049343e-21, -4.155564e-21, 
    2.098907e-20, -3.202631e-20, 2.152175e-20, 3.112696e-20, 2.617126e-20, 
    -1.740463e-20, 2.818826e-20, 1.259339e-20, 2.74475e-20, -5.271789e-21, 
    3.109983e-20, 2.119351e-20, 3.61149e-20, 2.296256e-20, -1.657623e-20, 
    -2.419035e-21, 3.408598e-21, -5.889198e-20, -2.173945e-20, -1.983158e-20, 
    7.406967e-21, -2.900678e-20, -4.06106e-20, 2.067497e-20, 1.850219e-20, 
    1.436836e-21, -2.124608e-20, 9.485329e-21, -1.206469e-20, 1.717504e-20, 
    7.461198e-22, -4.018462e-21, 1.252187e-20, -9.85714e-21, 1.825053e-20, 
    -9.162734e-21, -2.866778e-20, -1.350805e-20, -9.955797e-21, 
    -1.764353e-20, 2.758435e-20, -3.529949e-20, 4.392362e-20, 2.14177e-20, 
    -4.222755e-20, -1.052322e-21, -2.139621e-20, 2.080475e-20, -7.345346e-22, 
    5.399022e-21, -1.52525e-20, 8.114926e-21, -2.435642e-20, 8.129362e-21, 
    -1.134512e-20, 3.067515e-20, -8.188724e-21, 2.820381e-20, 4.89295e-21, 
    -2.857617e-20, 3.503883e-20, 1.233893e-20, -1.056141e-20, 4.845183e-20, 
    -7.181355e-21, -3.071474e-20, 3.084504e-23, -2.204395e-20, -4.202779e-21, 
    -1.705405e-20, 5.824259e-21, 2.832687e-21, 1.276814e-20, -8.632038e-21, 
    -2.598747e-20, 3.849861e-20, -2.004165e-20, 3.388612e-20, -8.602359e-21, 
    -1.97852e-20, 1.425359e-20, 5.463487e-21, 1.680015e-20, 1.287951e-20, 
    -6.317629e-21, 2.841558e-20, -6.212431e-21, 1.247663e-20, 2.952163e-20, 
    3.379905e-20, -9.723687e-21, 4.389479e-20, 2.356615e-20, -2.002157e-20, 
    -1.366409e-20, -1.511751e-21, 8.69171e-21, 7.705805e-21, -7.792053e-21, 
    -1.61295e-20, 3.983607e-22, -3.172803e-21, -1.726057e-21, 2.477683e-20, 
    2.203604e-20, -5.256824e-21, -4.188932e-21, -1.514419e-20, 2.148189e-20, 
    6.747096e-21, -3.566649e-21, -3.387567e-20, -2.46284e-20, -2.642289e-20, 
    -1.329004e-20, -9.560523e-21, -3.991141e-20, 1.356683e-20, -7.313102e-21, 
    -3.113147e-21, 7.868969e-21, -4.408961e-20, -6.698746e-21, -9.067112e-22, 
    -4.49881e-21, -1.566499e-20, 7.274808e-22, 2.540902e-20, 1.014807e-20, 
    -3.29449e-20, -1.831417e-20, -2.645369e-20, -3.638169e-21, -3.733147e-20, 
    2.509546e-20, 6.605454e-21, 2.253935e-21, -4.409215e-20, 8.001842e-23, 
    -1.316395e-20, 4.810664e-20, -1.5447e-20, -1.741733e-20, -4.415013e-20, 
    -2.137671e-20, 5.831902e-21, -1.455442e-20, -2.02017e-20, 3.93984e-21, 
    -1.48609e-20, -8.243849e-21, -1.039063e-20, 2.541466e-21, -3.108849e-20, 
    3.486338e-21, 8.535366e-21, -6.036286e-21, 2.993851e-21, 1.604792e-21, 
    2.996919e-20, -3.522797e-20, -1.5961e-20, 1.876492e-21, -6.754243e-22, 
    1.163662e-20, 2.46264e-20, 6.164654e-21, 6.123327e-20, 5.748226e-21, 
    -2.01932e-20, -2.4599e-20, 1.534946e-20, -1.992093e-20, 3.098305e-20, 
    2.824933e-20, 3.949467e-20, 1.126144e-20, 3.999172e-20, -1.13166e-20, 
    -4.343876e-21, -1.679223e-20, 7.08749e-21, -9.251807e-21, -2.195293e-20, 
    -1.471338e-21, -2.829767e-20, -7.141488e-21, -1.583717e-20, 4.489888e-22, 
    3.486917e-20, 1.148228e-20, 1.115852e-20, 1.703743e-21, -3.41239e-20, 
    4.367339e-21, 2.500724e-20, 1.86362e-20, -1.095158e-20, 3.742873e-20, 
    -2.430553e-20, 1.161601e-20, -2.044229e-20, -2.311211e-20, 2.219749e-20, 
    2.532392e-20, -2.706442e-20, -1.532145e-20, -6.36201e-21, -3.685762e-20, 
    2.294812e-20, 1.149498e-20, 4.040703e-20, -2.292976e-20, 1.989801e-20, 
    1.388576e-20, -8.291071e-21, 5.242961e-21, 4.987739e-20, -2.018615e-20, 
    -4.044466e-21, 3.38143e-20, 1.197056e-20, 1.690844e-20 ;

 M_SOIL2C_TO_LEACHING =
  1.002504e-20, 2.114231e-20, 1.763079e-20, 1.182013e-20, 1.225893e-20, 
    1.363038e-21, 6.741421e-21, -4.061726e-21, -3.490279e-21, 1.688892e-20, 
    -2.46612e-20, 2.513108e-20, -2.424274e-20, -3.733121e-20, -1.113309e-20, 
    -2.905852e-20, -2.317741e-20, 4.636192e-20, -4.32308e-22, -1.503226e-20, 
    1.971707e-20, 4.398463e-21, 4.403416e-20, -4.18679e-20, 1.257558e-20, 
    -1.164343e-20, -2.994994e-20, -3.02325e-21, 2.328203e-20, 1.469012e-20, 
    -1.531215e-20, 3.563708e-20, -1.840181e-20, 5.44511e-21, 6.822583e-21, 
    5.920664e-21, -1.395106e-20, 3.811178e-22, 9.896436e-21, -5.378726e-20, 
    2.046065e-20, 5.155578e-21, -2.588878e-20, -2.67384e-20, 3.53725e-21, 
    -1.446309e-20, 1.402432e-20, 9.96513e-21, 2.123021e-21, -2.373158e-20, 
    2.73203e-21, 1.046835e-20, 4.128548e-20, -1.212548e-20, 8.626673e-21, 
    -1.201437e-20, -4.223743e-20, -1.909196e-20, -8.758437e-21, 2.732536e-20, 
    -2.542894e-21, 5.800224e-21, -8.839289e-21, -3.408292e-20, -2.738672e-20, 
    -1.557822e-21, 3.867418e-20, 7.935123e-21, 1.559712e-20, 4.027923e-20, 
    1.325723e-20, 9.356978e-21, 2.343073e-20, 1.871535e-20, 2.827733e-20, 
    3.421072e-20, 9.854022e-21, -3.133135e-20, 3.453835e-21, 2.852383e-20, 
    -6.39264e-22, 1.286087e-20, 1.535961e-20, 2.538442e-20, 2.425604e-20, 
    -1.822509e-20, 3.590399e-20, 3.123102e-20, -6.088032e-21, 1.499208e-20, 
    3.171901e-20, -2.646473e-20, 1.982877e-20, 1.787254e-20, 3.07775e-20, 
    7.667099e-21, -2.561682e-20, 2.06747e-20, 2.524617e-20, -2.301824e-20, 
    1.40373e-20, 1.547398e-21, -6.237038e-21, -2.578504e-20, -1.810751e-20, 
    -1.055322e-20, -2.27946e-20, -4.1994e-21, 1.170249e-20, 2.955952e-21, 
    9.950433e-21, -2.191786e-20, 1.433021e-20, 1.386115e-20, 1.201889e-20, 
    -2.485483e-21, 8.353577e-21, -2.35198e-20, 2.169681e-21, -1.366691e-20, 
    4.48977e-21, 4.133948e-20, 9.027313e-21, 4.867664e-20, -2.919137e-20, 
    2.64636e-20, -1.117577e-20, 1.897801e-20, 3.230198e-20, -2.191475e-20, 
    2.139678e-20, 3.421946e-20, 4.937441e-20, 2.476835e-20, -4.076707e-21, 
    -5.510147e-21, 2.594109e-20, -3.077299e-20, 2.873111e-20, 2.723037e-20, 
    2.151616e-22, 1.078343e-21, -1.865089e-20, -4.24381e-22, -1.759154e-20, 
    -7.403503e-20, -1.832236e-20, -2.328287e-21, -2.550911e-20, 
    -2.948967e-20, 9.49921e-21, 2.392635e-20, -1.789686e-20, -1.363413e-20, 
    2.834603e-20, 9.066608e-21, -2.057235e-20, -6.686589e-21, 2.844287e-22, 
    -2.226503e-21, -3.359775e-20, 2.283022e-20, -3.038804e-21, 2.004336e-20, 
    2.715968e-20, 3.05058e-20, -8.752216e-21, -9.112678e-21, 1.303104e-21, 
    -3.143118e-20, -1.374077e-21, -3.785486e-21, -1.374525e-20, 1.882083e-20, 
    -3.038651e-20, 9.564492e-21, 5.723716e-20, 1.87846e-21, 2.662307e-20, 
    -1.573e-20, -4.736871e-20, 2.762365e-20, 1.630905e-20, -4.839078e-20, 
    1.506051e-20, 2.430778e-20, 2.372308e-20, -8.900404e-22, -5.575167e-21, 
    1.236071e-20, 3.318526e-20, 2.410986e-20, 4.415831e-20, -6.678401e-21, 
    -1.552051e-20, -1.931899e-20, 7.165523e-21, 2.865223e-20, 2.031335e-20, 
    -1.773175e-20, -1.623553e-20, -2.057235e-20, -6.004062e-21, 2.645372e-20, 
    -9.90971e-21, -1.994721e-20, 3.791334e-20, 2.955948e-20, -2.652409e-20, 
    2.344975e-21, -1.398074e-20, -1.633618e-20, 3.38177e-20, 9.280373e-21, 
    -3.041317e-21, 9.735272e-21, -1.63246e-20, 2.252912e-20, -1.226769e-20, 
    -4.301747e-21, -2.889565e-20, -9.844379e-21, -1.192846e-21, 
    -2.495892e-20, 2.949276e-20, 2.695641e-20, 1.178411e-21, -1.196714e-20, 
    -4.309651e-21, 1.059988e-20, 6.472262e-21, 5.523732e-21, -9.350185e-21, 
    -3.723845e-21, -1.861358e-20, 2.256134e-20, -1.938062e-20, -1.336356e-20, 
    -3.08742e-20, -2.117991e-20, -1.167136e-21, 1.37198e-20, 2.95403e-20, 
    -1.02241e-20, 1.954491e-20, 6.055807e-21, -2.997171e-20, 4.041279e-23, 
    4.914413e-21, -4.801337e-21, 6.935398e-21, 2.78491e-21, -2.157293e-20, 
    9.37818e-22, 2.230406e-20, -2.066173e-21, 1.202482e-20, 1.60263e-20, 
    1.297651e-20, 8.028988e-21, 6.191792e-21, 2.833923e-20, -4.685611e-20, 
    -1.788019e-20, -4.574869e-21, 2.904239e-20, -6.419205e-20, 8.219552e-21, 
    1.482412e-20, 1.284502e-20, 2.3854e-20, -3.496418e-20, 2.081491e-20, 
    2.329222e-20, 8.035138e-22, -6.581963e-21, -7.715993e-21, 8.068855e-21, 
    3.578807e-21, -2.429902e-20, -1.755558e-20, 7.478264e-22, -2.60087e-20, 
    7.307183e-21, -1.753779e-20, 5.736331e-21, 1.064479e-21, -8.816943e-21, 
    3.160081e-20, -2.43895e-20, 2.536376e-20, 3.147061e-21, 3.119351e-21, 
    -2.709013e-20, 2.703359e-20, -4.955452e-20, 2.948881e-21, 1.67826e-20, 
    -8.021633e-21, 5.202548e-21, 1.378622e-20, 5.366226e-21, -1.96865e-21, 
    2.999123e-20, 3.241e-20, 1.65679e-21, 4.088288e-20, 1.965545e-20, 
    -9.009791e-21, 4.472547e-20, -3.940814e-20, -4.391081e-21, -1.476955e-20, 
    1.781289e-20, -5.936217e-21, -2.345987e-20, 1.797745e-20, -9.843807e-21, 
    6.639646e-21, 2.182853e-20, -1.568816e-20, -4.239802e-20, -2.660355e-20, 
    -6.25487e-21, -4.469393e-21, -1.315261e-21, 1.193392e-21, -4.131065e-20, 
    8.637434e-21, 2.736893e-20, 3.891762e-20, -4.462877e-20, 1.057425e-21, 
    9.118144e-22, -5.346159e-21, 2.566487e-20, 1.771223e-20, 9.156798e-21 ;

 M_SOIL3C_TO_LEACHING =
  -1.288292e-20, 3.267066e-20, -1.757144e-20, -3.005697e-21, 2.941786e-20, 
    2.467392e-20, 1.33955e-20, 1.232649e-22, -1.291225e-21, -2.875289e-20, 
    2.006905e-20, 5.674707e-21, -7.11266e-21, -3.168289e-21, -4.704517e-22, 
    2.907179e-20, -2.626484e-20, 1.162758e-20, -2.976956e-20, 8.683522e-21, 
    3.350916e-21, 3.129557e-21, -2.189325e-20, -7.789202e-21, 1.291287e-20, 
    1.282437e-20, -1.104656e-20, -4.489486e-21, 1.360245e-20, 2.065066e-20, 
    2.929289e-20, 6.161551e-21, 1.397369e-20, -1.400845e-20, 1.169884e-20, 
    2.862534e-20, -1.162858e-21, -7.97046e-21, -3.961991e-20, 2.27714e-20, 
    -1.155634e-20, -2.68436e-20, 7.553712e-21, 3.011903e-20, 1.977021e-20, 
    3.549979e-21, -3.272059e-21, 2.992144e-21, -5.47282e-21, 4.002364e-21, 
    1.405566e-20, 1.95446e-20, 7.490364e-21, 3.024647e-21, -4.283369e-21, 
    1.559429e-20, 2.57025e-20, -3.771826e-20, -7.052987e-21, -1.53438e-20, 
    -2.408612e-20, -1.402401e-20, -1.86037e-20, -2.6195e-20, 1.447582e-20, 
    -2.849558e-20, -5.579269e-20, -5.034592e-21, 2.810324e-22, 6.009458e-21, 
    3.675496e-21, 1.12702e-20, 1.606023e-20, -4.018649e-20, -2.105809e-20, 
    3.066357e-20, 3.329071e-20, 1.40014e-20, 2.167159e-20, 1.961983e-20, 
    -2.791391e-21, -2.305982e-20, -1.932268e-20, 1.960426e-20, -8.44856e-21, 
    1.97004e-20, -2.960388e-20, -1.251678e-20, 2.123222e-20, -1.312715e-21, 
    4.665157e-22, 5.449069e-20, -3.683219e-20, -2.134364e-20, 2.193916e-22, 
    -2.252262e-20, -2.552635e-20, -2.302418e-20, 9.689184e-21, -3.954895e-20, 
    2.894427e-20, 9.194697e-21, -8.101652e-21, 2.754588e-20, -5.040812e-21, 
    6.378109e-21, 1.934925e-20, -1.927601e-20, 1.898311e-20, 1.043672e-20, 
    -2.841558e-20, 9.7073e-21, 1.779394e-20, 1.538704e-20, -2.908931e-20, 
    -3.537783e-20, -1.412635e-20, -2.05189e-20, 9.081076e-22, 8.883408e-21, 
    3.887549e-21, 8.108444e-21, -2.379603e-20, 2.880349e-20, -1.102255e-20, 
    -6.397058e-21, 6.352939e-21, -1.561218e-21, 3.61149e-20, 2.670704e-20, 
    -9.598421e-21, -1.038923e-20, 6.053546e-21, 1.867973e-20, -8.840717e-21, 
    2.031817e-20, -1.564319e-20, 1.378199e-20, 1.316847e-20, 2.010224e-21, 
    4.466948e-20, 4.212575e-20, -3.101562e-21, 1.802862e-20, 7.570409e-21, 
    -1.013788e-20, -2.516786e-20, 9.552351e-21, 1.764296e-20, 1.813423e-21, 
    6.849705e-21, 1.332963e-20, 3.610753e-20, -5.295376e-20, 2.26535e-20, 
    -1.595338e-20, 2.097071e-20, -4.156202e-22, -6.849704e-21, -7.589904e-21, 
    -1.051815e-20, 6.9775e-21, -1.705008e-20, 3.316149e-20, 1.687225e-20, 
    1.928734e-20, -1.751802e-20, 1.285315e-21, 2.33414e-20, 1.437008e-20, 
    -2.605761e-20, 4.268934e-21, -3.605683e-21, 1.586599e-20, 3.237353e-20, 
    -3.278999e-20, -2.070777e-20, 1.221455e-20, -1.420101e-20, -5.496855e-21, 
    5.117371e-23, -3.384284e-21, 1.119245e-20, 6.740849e-21, -5.417399e-21, 
    -1.929976e-20, 1.011186e-20, -3.453245e-20, 3.316177e-20, 1.077657e-20, 
    7.347033e-21, -2.262864e-20, 1.105818e-20, -3.969145e-20, -1.664296e-20, 
    -1.714395e-20, 4.827913e-21, -3.822858e-20, 2.474461e-20, 1.013931e-20, 
    5.342484e-21, 1.459654e-20, -1.4754e-20, -2.049883e-20, 8.503409e-21, 
    -3.135667e-22, -1.635425e-20, 8.351316e-21, -3.579768e-20, 1.264402e-20, 
    -7.814399e-21, -1.783013e-20, 9.27527e-21, -1.082859e-20, 1.085035e-20, 
    -1.968088e-20, 1.639329e-20, 1.488097e-20, 3.082585e-20, -2.700097e-22, 
    -1.500763e-20, 1.487021e-20, 1.088768e-20, 2.049629e-20, -1.691126e-20, 
    1.521431e-20, 3.394776e-20, -6.069438e-20, -2.632309e-20, 1.054499e-22, 
    1.918696e-20, 2.576802e-21, 2.022682e-20, 3.148768e-21, 2.80274e-20, 
    -2.13869e-20, -1.528727e-20, -4.795229e-22, -3.896737e-20, -1.60676e-21, 
    2.370105e-20, -2.798499e-20, -6.566721e-21, -4.052947e-20, 7.460991e-21, 
    1.16536e-20, -1.102707e-20, 2.591935e-20, -2.056752e-20, -1.216789e-20, 
    1.124474e-20, 2.734091e-20, 3.562047e-23, 8.07e-21, -4.167112e-20, 
    3.730638e-21, -2.362046e-20, 2.019206e-20, 3.398169e-20, -1.428722e-20, 
    2.503552e-20, -2.963896e-20, -3.628003e-20, 1.62412e-20, -2.627249e-20, 
    7.725327e-21, -8.999602e-21, -1.591774e-20, -5.118417e-20, -2.599511e-20, 
    8.162158e-21, 2.758095e-20, -1.069147e-20, -2.234421e-20, 3.729924e-20, 
    1.206554e-20, -3.958768e-20, -1.044323e-20, -1.693954e-20, 7.505111e-21, 
    -2.179828e-20, -1.840406e-20, -1.236468e-20, -1.025972e-20, 1.641224e-20, 
    2.076348e-20, -1.182946e-20, 1.348571e-20, 1.476875e-20, -1.722112e-20, 
    -1.510927e-21, 3.58271e-20, 1.47232e-20, 6.329786e-21, 1.261405e-20, 
    1.058602e-20, -2.343047e-20, -1.745013e-20, 2.030291e-21, -4.248455e-20, 
    1.907809e-20, -2.118953e-20, -9.306376e-21, -3.060872e-20, 5.304585e-21, 
    8.928649e-22, -3.503319e-21, -4.290977e-20, 1.068014e-20, -1.150123e-20, 
    1.340115e-20, 1.413597e-20, 2.17787e-21, -9.781931e-21, 1.644307e-20, 
    -1.689571e-20, 9.651874e-21, 4.348825e-20, 6.326935e-21, -6.522601e-21, 
    -2.807517e-21, 7.836173e-21, 6.639384e-21, 6.166303e-20, -7.337154e-21, 
    -1.130633e-21, -2.11952e-20, -2.653032e-20, -1.756719e-20, 4.43288e-20, 
    9.569594e-21, -1.636532e-20, -2.785605e-20, -3.762948e-20, -2.672428e-20, 
    4.588239e-20, -3.733657e-20, 1.555338e-23 ;

 NBP =
  -6.35757e-08, -6.385525e-08, -6.38009e-08, -6.402639e-08, -6.39013e-08, 
    -6.404895e-08, -6.363237e-08, -6.386636e-08, -6.371699e-08, 
    -6.360087e-08, -6.446398e-08, -6.403645e-08, -6.490803e-08, 
    -6.463537e-08, -6.532027e-08, -6.48656e-08, -6.541195e-08, -6.530715e-08, 
    -6.562256e-08, -6.55322e-08, -6.593564e-08, -6.566426e-08, -6.614476e-08, 
    -6.587083e-08, -6.591368e-08, -6.565531e-08, -6.412248e-08, 
    -6.441076e-08, -6.41054e-08, -6.41465e-08, -6.412806e-08, -6.390389e-08, 
    -6.379094e-08, -6.355432e-08, -6.359728e-08, -6.377105e-08, 
    -6.416499e-08, -6.403126e-08, -6.436827e-08, -6.436066e-08, 
    -6.473585e-08, -6.456669e-08, -6.519728e-08, -6.501806e-08, 
    -6.553597e-08, -6.540572e-08, -6.552985e-08, -6.549221e-08, 
    -6.553034e-08, -6.533932e-08, -6.542116e-08, -6.525307e-08, 
    -6.459837e-08, -6.479079e-08, -6.421691e-08, -6.387185e-08, 
    -6.364264e-08, -6.347999e-08, -6.350298e-08, -6.354682e-08, 
    -6.377208e-08, -6.398385e-08, -6.414524e-08, -6.42532e-08, -6.435957e-08, 
    -6.468156e-08, -6.485197e-08, -6.523354e-08, -6.516466e-08, 
    -6.528133e-08, -6.539276e-08, -6.557987e-08, -6.554907e-08, 
    -6.563151e-08, -6.527824e-08, -6.551303e-08, -6.512544e-08, 
    -6.523145e-08, -6.438852e-08, -6.406734e-08, -6.393085e-08, 
    -6.381136e-08, -6.352067e-08, -6.372141e-08, -6.364228e-08, 
    -6.383054e-08, -6.395017e-08, -6.3891e-08, -6.425615e-08, -6.411419e-08, 
    -6.486207e-08, -6.453993e-08, -6.537977e-08, -6.51788e-08, -6.542793e-08, 
    -6.53008e-08, -6.551863e-08, -6.532259e-08, -6.566219e-08, -6.573613e-08, 
    -6.56856e-08, -6.587971e-08, -6.531172e-08, -6.552985e-08, -6.388935e-08, 
    -6.389899e-08, -6.394394e-08, -6.374634e-08, -6.373425e-08, 
    -6.355315e-08, -6.371429e-08, -6.378291e-08, -6.39571e-08, -6.406013e-08, 
    -6.415808e-08, -6.437342e-08, -6.461393e-08, -6.495023e-08, 
    -6.519183e-08, -6.535377e-08, -6.525447e-08, -6.534214e-08, 
    -6.524414e-08, -6.519819e-08, -6.570843e-08, -6.542193e-08, 
    -6.585179e-08, -6.5828e-08, -6.563347e-08, -6.583068e-08, -6.390577e-08, 
    -6.385024e-08, -6.365745e-08, -6.380832e-08, -6.353343e-08, -6.36873e-08, 
    -6.377579e-08, -6.411717e-08, -6.419216e-08, -6.426171e-08, 
    -6.439907e-08, -6.457535e-08, -6.488458e-08, -6.515364e-08, 
    -6.539925e-08, -6.538125e-08, -6.538759e-08, -6.544246e-08, 
    -6.530654e-08, -6.546477e-08, -6.549133e-08, -6.542189e-08, 
    -6.582482e-08, -6.570971e-08, -6.58275e-08, -6.575254e-08, -6.386828e-08, 
    -6.396172e-08, -6.391124e-08, -6.400618e-08, -6.393929e-08, 
    -6.423671e-08, -6.432588e-08, -6.474312e-08, -6.457188e-08, 
    -6.484441e-08, -6.459956e-08, -6.464295e-08, -6.485331e-08, 
    -6.461279e-08, -6.513881e-08, -6.47822e-08, -6.544459e-08, -6.508849e-08, 
    -6.546691e-08, -6.539818e-08, -6.551196e-08, -6.561386e-08, 
    -6.574206e-08, -6.59786e-08, -6.592382e-08, -6.612164e-08, -6.410102e-08, 
    -6.422221e-08, -6.421153e-08, -6.433836e-08, -6.443215e-08, 
    -6.463544e-08, -6.496149e-08, -6.483888e-08, -6.506396e-08, 
    -6.510916e-08, -6.476719e-08, -6.497716e-08, -6.430331e-08, 
    -6.441219e-08, -6.434736e-08, -6.411058e-08, -6.486714e-08, 
    -6.447888e-08, -6.519582e-08, -6.498549e-08, -6.559934e-08, 
    -6.529407e-08, -6.589367e-08, -6.615002e-08, -6.639124e-08, 
    -6.667317e-08, -6.428834e-08, -6.4206e-08, -6.435344e-08, -6.455743e-08, 
    -6.47467e-08, -6.499832e-08, -6.502406e-08, -6.507121e-08, -6.51933e-08, 
    -6.529596e-08, -6.508611e-08, -6.53217e-08, -6.443745e-08, -6.490084e-08, 
    -6.417487e-08, -6.439348e-08, -6.454541e-08, -6.447876e-08, 
    -6.482487e-08, -6.490644e-08, -6.523793e-08, -6.506657e-08, 
    -6.608675e-08, -6.56354e-08, -6.688783e-08, -6.653783e-08, -6.417723e-08, 
    -6.428806e-08, -6.467379e-08, -6.449026e-08, -6.501512e-08, 
    -6.514431e-08, -6.524932e-08, -6.538358e-08, -6.539807e-08, 
    -6.547761e-08, -6.534727e-08, -6.547247e-08, -6.499886e-08, -6.52105e-08, 
    -6.46297e-08, -6.477106e-08, -6.470603e-08, -6.463469e-08, -6.485485e-08, 
    -6.508942e-08, -6.509442e-08, -6.516963e-08, -6.53816e-08, -6.501724e-08, 
    -6.614502e-08, -6.544855e-08, -6.440892e-08, -6.462241e-08, 
    -6.465289e-08, -6.457019e-08, -6.513136e-08, -6.492802e-08, 
    -6.547567e-08, -6.532767e-08, -6.557018e-08, -6.544967e-08, 
    -6.543194e-08, -6.527716e-08, -6.51808e-08, -6.493735e-08, -6.473926e-08, 
    -6.458218e-08, -6.46187e-08, -6.479126e-08, -6.510376e-08, -6.539939e-08, 
    -6.533463e-08, -6.555175e-08, -6.497706e-08, -6.521804e-08, 
    -6.512491e-08, -6.536776e-08, -6.483562e-08, -6.528879e-08, 
    -6.471979e-08, -6.476968e-08, -6.492399e-08, -6.52344e-08, -6.530306e-08, 
    -6.537638e-08, -6.533113e-08, -6.51117e-08, -6.507574e-08, -6.492024e-08, 
    -6.487731e-08, -6.475882e-08, -6.466072e-08, -6.475035e-08, 
    -6.484448e-08, -6.511178e-08, -6.535268e-08, -6.561532e-08, 
    -6.567959e-08, -6.598647e-08, -6.573666e-08, -6.61489e-08, -6.579844e-08, 
    -6.64051e-08, -6.531504e-08, -6.578811e-08, -6.493101e-08, -6.502334e-08, 
    -6.519036e-08, -6.557342e-08, -6.536661e-08, -6.560847e-08, 
    -6.507433e-08, -6.479721e-08, -6.47255e-08, -6.459173e-08, -6.472857e-08, 
    -6.471743e-08, -6.484837e-08, -6.480629e-08, -6.512066e-08, -6.49518e-08, 
    -6.54315e-08, -6.560656e-08, -6.610091e-08, -6.640397e-08, -6.671245e-08, 
    -6.684864e-08, -6.689009e-08, -6.690742e-08 ;

 NDEPLOY =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NDEP_TO_SMINN =
  3.989144e-10, 3.989147e-10, 3.989121e-10, 3.989123e-10, 3.989108e-10, 
    3.989089e-10, 3.989084e-10, 3.989066e-10, 3.98906e-10, 3.989042e-10, 
    3.989026e-10, 3.989029e-10, 3.989014e-10, 3.988995e-10, 3.988979e-10, 
    3.988982e-10, 3.988966e-10, 3.988948e-10, 3.988943e-10, 3.988924e-10, 
    3.988909e-10, 3.988911e-10, 3.988885e-10, 3.988888e-10, 3.988872e-10, 
    3.988854e-10, 3.989112e-10, 3.989115e-10, 3.989089e-10, 3.989092e-10, 
    3.989076e-10, 3.989057e-10, 3.989052e-10, 3.989034e-10, 3.989018e-10, 
    3.989021e-10, 3.989005e-10, 3.988987e-10, 3.988971e-10, 3.988974e-10, 
    3.988947e-10, 3.98895e-10, 3.988934e-10, 3.988916e-10, 3.988911e-10, 
    3.988892e-10, 3.988887e-10, 3.988869e-10, 3.988853e-10, 3.988856e-10, 
    3.98883e-10, 3.988832e-10, 3.989091e-10, 3.989072e-10, 3.989067e-10, 
    3.989049e-10, 3.989033e-10, 3.989036e-10, 3.98901e-10, 3.989012e-10, 
    3.988997e-10, 3.988978e-10, 3.988973e-10, 3.988955e-10, 3.988939e-10, 
    3.988942e-10, 3.988926e-10, 3.988908e-10, 3.988903e-10, 3.988884e-10, 
    3.988879e-10, 3.98886e-10, 3.988855e-10, 3.988837e-10, 3.988821e-10, 
    3.988824e-10, 3.988798e-10, 3.9888e-10, 3.989059e-10, 3.98904e-10, 
    3.989035e-10, 3.989017e-10, 3.989001e-10, 3.989004e-10, 3.988988e-10, 
    3.98897e-10, 3.988965e-10, 3.988946e-10, 3.988941e-10, 3.988923e-10, 
    3.988907e-10, 3.98891e-10, 3.988894e-10, 3.988876e-10, 3.98886e-10, 
    3.988863e-10, 3.988836e-10, 3.988839e-10, 3.988813e-10, 3.988816e-10, 
    3.988789e-10, 3.988792e-10, 3.988766e-10, 3.988768e-10, 3.989017e-10, 
    3.989019e-10, 3.989004e-10, 3.988985e-10, 3.98898e-10, 3.988962e-10, 
    3.988946e-10, 3.988949e-10, 3.988933e-10, 3.988914e-10, 3.988899e-10, 
    3.988901e-10, 3.988886e-10, 3.988867e-10, 3.988862e-10, 3.988844e-10, 
    3.988839e-10, 3.98882e-10, 3.988815e-10, 3.988797e-10, 3.988781e-10, 
    3.988784e-10, 3.988757e-10, 3.98876e-10, 3.988744e-10, 3.988726e-10, 
    3.988995e-10, 3.988977e-10, 3.988972e-10, 3.988953e-10, 3.988938e-10, 
    3.98894e-10, 3.988924e-10, 3.988906e-10, 3.98889e-10, 3.988893e-10, 
    3.988878e-10, 3.988859e-10, 3.988854e-10, 3.988835e-10, 3.98883e-10, 
    3.988812e-10, 3.988807e-10, 3.988788e-10, 3.988783e-10, 3.988765e-10, 
    3.988749e-10, 3.988752e-10, 3.988725e-10, 3.988728e-10, 3.988712e-10, 
    3.988694e-10, 3.988963e-10, 3.988945e-10, 3.988929e-10, 3.988932e-10, 
    3.988906e-10, 3.988908e-10, 3.988893e-10, 3.988874e-10, 3.988858e-10, 
    3.988861e-10, 3.988835e-10, 3.988838e-10, 3.988822e-10, 3.988803e-10, 
    3.988798e-10, 3.98878e-10, 3.988775e-10, 3.988756e-10, 3.988751e-10, 
    3.988733e-10, 3.988717e-10, 3.98872e-10, 3.988694e-10, 3.988696e-10, 
    3.98867e-10, 3.988673e-10, 3.988931e-10, 3.988913e-10, 3.988908e-10, 
    3.988889e-10, 3.988874e-10, 3.988876e-10, 3.988861e-10, 3.988842e-10, 
    3.988826e-10, 3.988829e-10, 3.988803e-10, 3.988806e-10, 3.98879e-10, 
    3.988772e-10, 3.988767e-10, 3.988748e-10, 3.988743e-10, 3.988724e-10, 
    3.988719e-10, 3.988701e-10, 3.988685e-10, 3.988688e-10, 3.988662e-10, 
    3.988664e-10, 3.988649e-10, 3.98863e-10, 3.988899e-10, 3.988881e-10, 
    3.988865e-10, 3.988868e-10, 3.988842e-10, 3.988845e-10, 3.988829e-10, 
    3.98881e-10, 3.988795e-10, 3.988797e-10, 3.988782e-10, 3.988763e-10, 
    3.988758e-10, 3.98874e-10, 3.988724e-10, 3.988727e-10, 3.9887e-10, 
    3.988703e-10, 3.988687e-10, 3.988669e-10, 3.988653e-10, 3.988656e-10, 
    3.98863e-10, 3.988632e-10, 3.988606e-10, 3.988609e-10, 3.988868e-10, 
    3.988849e-10, 3.988833e-10, 3.988836e-10, 3.98881e-10, 3.988813e-10, 
    3.988786e-10, 3.988789e-10, 3.988763e-10, 3.988765e-10, 3.988739e-10, 
    3.988742e-10, 3.988716e-10, 3.988719e-10, 3.988703e-10, 3.988684e-10, 
    3.988679e-10, 3.988661e-10, 3.988645e-10, 3.988648e-10, 3.988632e-10, 
    3.988614e-10, 3.988609e-10, 3.98859e-10, 3.988585e-10, 3.988566e-10, 
    3.988836e-10, 3.988817e-10, 3.988802e-10, 3.988804e-10, 3.988778e-10, 
    3.988781e-10, 3.988765e-10, 3.988747e-10, 3.988731e-10, 3.988734e-10, 
    3.988707e-10, 3.98871e-10, 3.988684e-10, 3.988687e-10, 3.98866e-10, 
    3.988663e-10, 3.988637e-10, 3.988639e-10, 3.988613e-10, 3.988616e-10, 
    3.9886e-10, 3.988582e-10, 3.988566e-10, 3.988569e-10, 3.988542e-10, 
    3.988545e-10, 3.988793e-10, 3.988796e-10, 3.98878e-10, 3.988762e-10, 
    3.988746e-10, 3.988749e-10, 3.988722e-10, 3.988725e-10, 3.988699e-10, 
    3.988702e-10, 3.988686e-10, 3.988667e-10, 3.988652e-10, 3.988655e-10, 
    3.988628e-10, 3.988631e-10, 3.988605e-10, 3.988607e-10, 3.988592e-10, 
    3.988573e-10, 3.988568e-10, 3.98855e-10, 3.988545e-10, 3.988526e-10, 
    3.988521e-10, 3.988503e-10, 3.988761e-10, 3.988764e-10, 3.988748e-10, 
    3.98873e-10, 3.988725e-10, 3.988706e-10, 3.98869e-10, 3.988693e-10, 
    3.988678e-10, 3.988659e-10, 3.988644e-10, 3.988646e-10, 3.98862e-10, 
    3.988623e-10, 3.988607e-10, 3.988589e-10, 3.988573e-10, 3.988576e-10, 
    3.988549e-10, 3.988552e-10, 3.988536e-10, 3.988518e-10, 3.988513e-10, 
    3.988494e-10, 3.988489e-10, 3.988476e-10 ;

 NEE =
  6.35757e-08, 6.385525e-08, 6.38009e-08, 6.402639e-08, 6.39013e-08, 
    6.404895e-08, 6.363237e-08, 6.386636e-08, 6.371699e-08, 6.360087e-08, 
    6.446398e-08, 6.403645e-08, 6.490803e-08, 6.463537e-08, 6.532027e-08, 
    6.48656e-08, 6.541195e-08, 6.530715e-08, 6.562256e-08, 6.55322e-08, 
    6.593564e-08, 6.566426e-08, 6.614476e-08, 6.587083e-08, 6.591368e-08, 
    6.565531e-08, 6.412248e-08, 6.441076e-08, 6.41054e-08, 6.41465e-08, 
    6.412806e-08, 6.390389e-08, 6.379094e-08, 6.355432e-08, 6.359728e-08, 
    6.377105e-08, 6.416499e-08, 6.403126e-08, 6.436827e-08, 6.436066e-08, 
    6.473585e-08, 6.456669e-08, 6.519728e-08, 6.501806e-08, 6.553597e-08, 
    6.540572e-08, 6.552985e-08, 6.549221e-08, 6.553034e-08, 6.533932e-08, 
    6.542116e-08, 6.525307e-08, 6.459837e-08, 6.479079e-08, 6.421691e-08, 
    6.387185e-08, 6.364264e-08, 6.347999e-08, 6.350298e-08, 6.354682e-08, 
    6.377208e-08, 6.398385e-08, 6.414524e-08, 6.42532e-08, 6.435957e-08, 
    6.468156e-08, 6.485197e-08, 6.523354e-08, 6.516466e-08, 6.528133e-08, 
    6.539276e-08, 6.557987e-08, 6.554907e-08, 6.563151e-08, 6.527824e-08, 
    6.551303e-08, 6.512544e-08, 6.523145e-08, 6.438852e-08, 6.406734e-08, 
    6.393085e-08, 6.381136e-08, 6.352067e-08, 6.372141e-08, 6.364228e-08, 
    6.383054e-08, 6.395017e-08, 6.3891e-08, 6.425615e-08, 6.411419e-08, 
    6.486207e-08, 6.453993e-08, 6.537977e-08, 6.51788e-08, 6.542793e-08, 
    6.53008e-08, 6.551863e-08, 6.532259e-08, 6.566219e-08, 6.573613e-08, 
    6.56856e-08, 6.587971e-08, 6.531172e-08, 6.552985e-08, 6.388935e-08, 
    6.389899e-08, 6.394394e-08, 6.374634e-08, 6.373425e-08, 6.355315e-08, 
    6.371429e-08, 6.378291e-08, 6.39571e-08, 6.406013e-08, 6.415808e-08, 
    6.437342e-08, 6.461393e-08, 6.495023e-08, 6.519183e-08, 6.535377e-08, 
    6.525447e-08, 6.534214e-08, 6.524414e-08, 6.519819e-08, 6.570843e-08, 
    6.542193e-08, 6.585179e-08, 6.5828e-08, 6.563347e-08, 6.583068e-08, 
    6.390577e-08, 6.385024e-08, 6.365745e-08, 6.380832e-08, 6.353343e-08, 
    6.36873e-08, 6.377579e-08, 6.411717e-08, 6.419216e-08, 6.426171e-08, 
    6.439907e-08, 6.457535e-08, 6.488458e-08, 6.515364e-08, 6.539925e-08, 
    6.538125e-08, 6.538759e-08, 6.544246e-08, 6.530654e-08, 6.546477e-08, 
    6.549133e-08, 6.542189e-08, 6.582482e-08, 6.570971e-08, 6.58275e-08, 
    6.575254e-08, 6.386828e-08, 6.396172e-08, 6.391124e-08, 6.400618e-08, 
    6.393929e-08, 6.423671e-08, 6.432588e-08, 6.474312e-08, 6.457188e-08, 
    6.484441e-08, 6.459956e-08, 6.464295e-08, 6.485331e-08, 6.461279e-08, 
    6.513881e-08, 6.47822e-08, 6.544459e-08, 6.508849e-08, 6.546691e-08, 
    6.539818e-08, 6.551196e-08, 6.561386e-08, 6.574206e-08, 6.59786e-08, 
    6.592382e-08, 6.612164e-08, 6.410102e-08, 6.422221e-08, 6.421153e-08, 
    6.433836e-08, 6.443215e-08, 6.463544e-08, 6.496149e-08, 6.483888e-08, 
    6.506396e-08, 6.510916e-08, 6.476719e-08, 6.497716e-08, 6.430331e-08, 
    6.441219e-08, 6.434736e-08, 6.411058e-08, 6.486714e-08, 6.447888e-08, 
    6.519582e-08, 6.498549e-08, 6.559934e-08, 6.529407e-08, 6.589367e-08, 
    6.615002e-08, 6.639124e-08, 6.667317e-08, 6.428834e-08, 6.4206e-08, 
    6.435344e-08, 6.455743e-08, 6.47467e-08, 6.499832e-08, 6.502406e-08, 
    6.507121e-08, 6.51933e-08, 6.529596e-08, 6.508611e-08, 6.53217e-08, 
    6.443745e-08, 6.490084e-08, 6.417487e-08, 6.439348e-08, 6.454541e-08, 
    6.447876e-08, 6.482487e-08, 6.490644e-08, 6.523793e-08, 6.506657e-08, 
    6.608675e-08, 6.56354e-08, 6.688783e-08, 6.653783e-08, 6.417723e-08, 
    6.428806e-08, 6.467379e-08, 6.449026e-08, 6.501512e-08, 6.514431e-08, 
    6.524932e-08, 6.538358e-08, 6.539807e-08, 6.547761e-08, 6.534727e-08, 
    6.547247e-08, 6.499886e-08, 6.52105e-08, 6.46297e-08, 6.477106e-08, 
    6.470603e-08, 6.463469e-08, 6.485485e-08, 6.508942e-08, 6.509442e-08, 
    6.516963e-08, 6.53816e-08, 6.501724e-08, 6.614502e-08, 6.544855e-08, 
    6.440892e-08, 6.462241e-08, 6.465289e-08, 6.457019e-08, 6.513136e-08, 
    6.492802e-08, 6.547567e-08, 6.532767e-08, 6.557018e-08, 6.544967e-08, 
    6.543194e-08, 6.527716e-08, 6.51808e-08, 6.493735e-08, 6.473926e-08, 
    6.458218e-08, 6.46187e-08, 6.479126e-08, 6.510376e-08, 6.539939e-08, 
    6.533463e-08, 6.555175e-08, 6.497706e-08, 6.521804e-08, 6.512491e-08, 
    6.536776e-08, 6.483562e-08, 6.528879e-08, 6.471979e-08, 6.476968e-08, 
    6.492399e-08, 6.52344e-08, 6.530306e-08, 6.537638e-08, 6.533113e-08, 
    6.51117e-08, 6.507574e-08, 6.492024e-08, 6.487731e-08, 6.475882e-08, 
    6.466072e-08, 6.475035e-08, 6.484448e-08, 6.511178e-08, 6.535268e-08, 
    6.561532e-08, 6.567959e-08, 6.598647e-08, 6.573666e-08, 6.61489e-08, 
    6.579844e-08, 6.64051e-08, 6.531504e-08, 6.578811e-08, 6.493101e-08, 
    6.502334e-08, 6.519036e-08, 6.557342e-08, 6.536661e-08, 6.560847e-08, 
    6.507433e-08, 6.479721e-08, 6.47255e-08, 6.459173e-08, 6.472857e-08, 
    6.471743e-08, 6.484837e-08, 6.480629e-08, 6.512066e-08, 6.49518e-08, 
    6.54315e-08, 6.560656e-08, 6.610091e-08, 6.640397e-08, 6.671245e-08, 
    6.684864e-08, 6.689009e-08, 6.690742e-08 ;

 NEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NEP =
  -6.35757e-08, -6.385525e-08, -6.38009e-08, -6.402639e-08, -6.39013e-08, 
    -6.404895e-08, -6.363237e-08, -6.386636e-08, -6.371699e-08, 
    -6.360087e-08, -6.446398e-08, -6.403645e-08, -6.490803e-08, 
    -6.463537e-08, -6.532027e-08, -6.48656e-08, -6.541195e-08, -6.530715e-08, 
    -6.562256e-08, -6.55322e-08, -6.593564e-08, -6.566426e-08, -6.614476e-08, 
    -6.587083e-08, -6.591368e-08, -6.565531e-08, -6.412248e-08, 
    -6.441076e-08, -6.41054e-08, -6.41465e-08, -6.412806e-08, -6.390389e-08, 
    -6.379094e-08, -6.355432e-08, -6.359728e-08, -6.377105e-08, 
    -6.416499e-08, -6.403126e-08, -6.436827e-08, -6.436066e-08, 
    -6.473585e-08, -6.456669e-08, -6.519728e-08, -6.501806e-08, 
    -6.553597e-08, -6.540572e-08, -6.552985e-08, -6.549221e-08, 
    -6.553034e-08, -6.533932e-08, -6.542116e-08, -6.525307e-08, 
    -6.459837e-08, -6.479079e-08, -6.421691e-08, -6.387185e-08, 
    -6.364264e-08, -6.347999e-08, -6.350298e-08, -6.354682e-08, 
    -6.377208e-08, -6.398385e-08, -6.414524e-08, -6.42532e-08, -6.435957e-08, 
    -6.468156e-08, -6.485197e-08, -6.523354e-08, -6.516466e-08, 
    -6.528133e-08, -6.539276e-08, -6.557987e-08, -6.554907e-08, 
    -6.563151e-08, -6.527824e-08, -6.551303e-08, -6.512544e-08, 
    -6.523145e-08, -6.438852e-08, -6.406734e-08, -6.393085e-08, 
    -6.381136e-08, -6.352067e-08, -6.372141e-08, -6.364228e-08, 
    -6.383054e-08, -6.395017e-08, -6.3891e-08, -6.425615e-08, -6.411419e-08, 
    -6.486207e-08, -6.453993e-08, -6.537977e-08, -6.51788e-08, -6.542793e-08, 
    -6.53008e-08, -6.551863e-08, -6.532259e-08, -6.566219e-08, -6.573613e-08, 
    -6.56856e-08, -6.587971e-08, -6.531172e-08, -6.552985e-08, -6.388935e-08, 
    -6.389899e-08, -6.394394e-08, -6.374634e-08, -6.373425e-08, 
    -6.355315e-08, -6.371429e-08, -6.378291e-08, -6.39571e-08, -6.406013e-08, 
    -6.415808e-08, -6.437342e-08, -6.461393e-08, -6.495023e-08, 
    -6.519183e-08, -6.535377e-08, -6.525447e-08, -6.534214e-08, 
    -6.524414e-08, -6.519819e-08, -6.570843e-08, -6.542193e-08, 
    -6.585179e-08, -6.5828e-08, -6.563347e-08, -6.583068e-08, -6.390577e-08, 
    -6.385024e-08, -6.365745e-08, -6.380832e-08, -6.353343e-08, -6.36873e-08, 
    -6.377579e-08, -6.411717e-08, -6.419216e-08, -6.426171e-08, 
    -6.439907e-08, -6.457535e-08, -6.488458e-08, -6.515364e-08, 
    -6.539925e-08, -6.538125e-08, -6.538759e-08, -6.544246e-08, 
    -6.530654e-08, -6.546477e-08, -6.549133e-08, -6.542189e-08, 
    -6.582482e-08, -6.570971e-08, -6.58275e-08, -6.575254e-08, -6.386828e-08, 
    -6.396172e-08, -6.391124e-08, -6.400618e-08, -6.393929e-08, 
    -6.423671e-08, -6.432588e-08, -6.474312e-08, -6.457188e-08, 
    -6.484441e-08, -6.459956e-08, -6.464295e-08, -6.485331e-08, 
    -6.461279e-08, -6.513881e-08, -6.47822e-08, -6.544459e-08, -6.508849e-08, 
    -6.546691e-08, -6.539818e-08, -6.551196e-08, -6.561386e-08, 
    -6.574206e-08, -6.59786e-08, -6.592382e-08, -6.612164e-08, -6.410102e-08, 
    -6.422221e-08, -6.421153e-08, -6.433836e-08, -6.443215e-08, 
    -6.463544e-08, -6.496149e-08, -6.483888e-08, -6.506396e-08, 
    -6.510916e-08, -6.476719e-08, -6.497716e-08, -6.430331e-08, 
    -6.441219e-08, -6.434736e-08, -6.411058e-08, -6.486714e-08, 
    -6.447888e-08, -6.519582e-08, -6.498549e-08, -6.559934e-08, 
    -6.529407e-08, -6.589367e-08, -6.615002e-08, -6.639124e-08, 
    -6.667317e-08, -6.428834e-08, -6.4206e-08, -6.435344e-08, -6.455743e-08, 
    -6.47467e-08, -6.499832e-08, -6.502406e-08, -6.507121e-08, -6.51933e-08, 
    -6.529596e-08, -6.508611e-08, -6.53217e-08, -6.443745e-08, -6.490084e-08, 
    -6.417487e-08, -6.439348e-08, -6.454541e-08, -6.447876e-08, 
    -6.482487e-08, -6.490644e-08, -6.523793e-08, -6.506657e-08, 
    -6.608675e-08, -6.56354e-08, -6.688783e-08, -6.653783e-08, -6.417723e-08, 
    -6.428806e-08, -6.467379e-08, -6.449026e-08, -6.501512e-08, 
    -6.514431e-08, -6.524932e-08, -6.538358e-08, -6.539807e-08, 
    -6.547761e-08, -6.534727e-08, -6.547247e-08, -6.499886e-08, -6.52105e-08, 
    -6.46297e-08, -6.477106e-08, -6.470603e-08, -6.463469e-08, -6.485485e-08, 
    -6.508942e-08, -6.509442e-08, -6.516963e-08, -6.53816e-08, -6.501724e-08, 
    -6.614502e-08, -6.544855e-08, -6.440892e-08, -6.462241e-08, 
    -6.465289e-08, -6.457019e-08, -6.513136e-08, -6.492802e-08, 
    -6.547567e-08, -6.532767e-08, -6.557018e-08, -6.544967e-08, 
    -6.543194e-08, -6.527716e-08, -6.51808e-08, -6.493735e-08, -6.473926e-08, 
    -6.458218e-08, -6.46187e-08, -6.479126e-08, -6.510376e-08, -6.539939e-08, 
    -6.533463e-08, -6.555175e-08, -6.497706e-08, -6.521804e-08, 
    -6.512491e-08, -6.536776e-08, -6.483562e-08, -6.528879e-08, 
    -6.471979e-08, -6.476968e-08, -6.492399e-08, -6.52344e-08, -6.530306e-08, 
    -6.537638e-08, -6.533113e-08, -6.51117e-08, -6.507574e-08, -6.492024e-08, 
    -6.487731e-08, -6.475882e-08, -6.466072e-08, -6.475035e-08, 
    -6.484448e-08, -6.511178e-08, -6.535268e-08, -6.561532e-08, 
    -6.567959e-08, -6.598647e-08, -6.573666e-08, -6.61489e-08, -6.579844e-08, 
    -6.64051e-08, -6.531504e-08, -6.578811e-08, -6.493101e-08, -6.502334e-08, 
    -6.519036e-08, -6.557342e-08, -6.536661e-08, -6.560847e-08, 
    -6.507433e-08, -6.479721e-08, -6.47255e-08, -6.459173e-08, -6.472857e-08, 
    -6.471743e-08, -6.484837e-08, -6.480629e-08, -6.512066e-08, -6.49518e-08, 
    -6.54315e-08, -6.560656e-08, -6.610091e-08, -6.640397e-08, -6.671245e-08, 
    -6.684864e-08, -6.689009e-08, -6.690742e-08 ;

 NET_NMIN =
  8.956404e-09, 8.995784e-09, 8.988128e-09, 9.019892e-09, 9.002271e-09, 
    9.02307e-09, 8.964387e-09, 8.997348e-09, 8.976306e-09, 8.959948e-09, 
    9.081533e-09, 9.021308e-09, 9.144085e-09, 9.105678e-09, 9.202157e-09, 
    9.138109e-09, 9.215071e-09, 9.200308e-09, 9.244739e-09, 9.232011e-09, 
    9.288842e-09, 9.250614e-09, 9.3183e-09, 9.279711e-09, 9.285748e-09, 
    9.249352e-09, 9.033427e-09, 9.074036e-09, 9.031021e-09, 9.036812e-09, 
    9.034213e-09, 9.002636e-09, 8.986723e-09, 8.953393e-09, 8.959444e-09, 
    8.983923e-09, 9.039416e-09, 9.020578e-09, 9.068052e-09, 9.06698e-09, 
    9.119832e-09, 9.096002e-09, 9.184832e-09, 9.159585e-09, 9.232542e-09, 
    9.214194e-09, 9.23168e-09, 9.226378e-09, 9.231749e-09, 9.20484e-09, 
    9.216369e-09, 9.192691e-09, 9.100465e-09, 9.127571e-09, 9.04673e-09, 
    8.998122e-09, 8.965833e-09, 8.942921e-09, 8.94616e-09, 8.952335e-09, 
    8.984067e-09, 9.013899e-09, 9.036634e-09, 9.051842e-09, 9.066826e-09, 
    9.112184e-09, 9.136189e-09, 9.189939e-09, 9.180237e-09, 9.196671e-09, 
    9.212369e-09, 9.238725e-09, 9.234387e-09, 9.246e-09, 9.196237e-09, 
    9.22931e-09, 9.174712e-09, 9.189645e-09, 9.070903e-09, 9.02566e-09, 
    9.006433e-09, 8.9896e-09, 8.948651e-09, 8.976929e-09, 8.965782e-09, 
    8.992302e-09, 9.009154e-09, 9.00082e-09, 9.052258e-09, 9.03226e-09, 
    9.137612e-09, 9.092234e-09, 9.210538e-09, 9.182228e-09, 9.217323e-09, 
    9.199415e-09, 9.2301e-09, 9.202483e-09, 9.250321e-09, 9.260738e-09, 
    9.253619e-09, 9.280963e-09, 9.200953e-09, 9.23168e-09, 9.000586e-09, 
    9.001945e-09, 9.008278e-09, 8.980441e-09, 8.978739e-09, 8.953227e-09, 
    8.975927e-09, 8.985593e-09, 9.01013e-09, 9.024645e-09, 9.038442e-09, 
    9.068778e-09, 9.102657e-09, 9.15003e-09, 9.184063e-09, 9.206877e-09, 
    9.192887e-09, 9.205238e-09, 9.191432e-09, 9.18496e-09, 9.256835e-09, 
    9.216477e-09, 9.27703e-09, 9.27368e-09, 9.246276e-09, 9.274057e-09, 
    9.0029e-09, 8.995078e-09, 8.967919e-09, 8.989173e-09, 8.950449e-09, 
    8.972125e-09, 8.984589e-09, 9.032679e-09, 9.043243e-09, 9.053041e-09, 
    9.07239e-09, 9.097222e-09, 9.140783e-09, 9.178684e-09, 9.213282e-09, 
    9.210747e-09, 9.211639e-09, 9.219368e-09, 9.200223e-09, 9.222512e-09, 
    9.226253e-09, 9.216472e-09, 9.27323e-09, 9.257015e-09, 9.273609e-09, 
    9.26305e-09, 8.99762e-09, 9.010782e-09, 9.00367e-09, 9.017044e-09, 
    9.007622e-09, 9.049519e-09, 9.06208e-09, 9.120856e-09, 9.096733e-09, 
    9.135124e-09, 9.100632e-09, 9.106745e-09, 9.136377e-09, 9.102497e-09, 
    9.176595e-09, 9.12636e-09, 9.219669e-09, 9.169507e-09, 9.222813e-09, 
    9.213132e-09, 9.22916e-09, 9.243514e-09, 9.261572e-09, 9.294893e-09, 
    9.287177e-09, 9.315042e-09, 9.030404e-09, 9.047476e-09, 9.045972e-09, 
    9.063838e-09, 9.07705e-09, 9.105687e-09, 9.151616e-09, 9.134345e-09, 
    9.166052e-09, 9.172417e-09, 9.124246e-09, 9.153823e-09, 9.058901e-09, 
    9.074238e-09, 9.065106e-09, 9.03175e-09, 9.138326e-09, 9.083633e-09, 
    9.184626e-09, 9.154998e-09, 9.241467e-09, 9.198465e-09, 9.28293e-09, 
    9.31904e-09, 9.35302e-09, 9.392735e-09, 9.056793e-09, 9.045192e-09, 
    9.065962e-09, 9.094698e-09, 9.12136e-09, 9.156805e-09, 9.160431e-09, 
    9.167072e-09, 9.184271e-09, 9.198732e-09, 9.169172e-09, 9.202358e-09, 
    9.077796e-09, 9.143073e-09, 9.040807e-09, 9.071603e-09, 9.093005e-09, 
    9.083616e-09, 9.13237e-09, 9.143862e-09, 9.190557e-09, 9.166418e-09, 
    9.310128e-09, 9.246548e-09, 9.422972e-09, 9.37367e-09, 9.041139e-09, 
    9.056752e-09, 9.11109e-09, 9.085236e-09, 9.15917e-09, 9.177369e-09, 
    9.192163e-09, 9.211075e-09, 9.213116e-09, 9.224322e-09, 9.20596e-09, 
    9.223596e-09, 9.156881e-09, 9.186694e-09, 9.104878e-09, 9.124792e-09, 
    9.11563e-09, 9.105582e-09, 9.136595e-09, 9.169637e-09, 9.170342e-09, 
    9.180937e-09, 9.210796e-09, 9.159471e-09, 9.318336e-09, 9.220227e-09, 
    9.073776e-09, 9.10385e-09, 9.108144e-09, 9.096495e-09, 9.175545e-09, 
    9.146903e-09, 9.224048e-09, 9.203198e-09, 9.23736e-09, 9.220384e-09, 
    9.217888e-09, 9.196084e-09, 9.182511e-09, 9.148216e-09, 9.120313e-09, 
    9.098184e-09, 9.10333e-09, 9.127636e-09, 9.171658e-09, 9.213302e-09, 
    9.20418e-09, 9.234764e-09, 9.15381e-09, 9.187756e-09, 9.174636e-09, 
    9.208846e-09, 9.133886e-09, 9.197723e-09, 9.117569e-09, 9.124596e-09, 
    9.146334e-09, 9.190059e-09, 9.199732e-09, 9.210061e-09, 9.203687e-09, 
    9.172775e-09, 9.167711e-09, 9.145806e-09, 9.139758e-09, 9.123067e-09, 
    9.109248e-09, 9.121874e-09, 9.135134e-09, 9.172788e-09, 9.206722e-09, 
    9.243719e-09, 9.252772e-09, 9.296001e-09, 9.260813e-09, 9.318883e-09, 
    9.269515e-09, 9.354972e-09, 9.201419e-09, 9.268061e-09, 9.147323e-09, 
    9.16033e-09, 9.183857e-09, 9.237817e-09, 9.208684e-09, 9.242754e-09, 
    9.167512e-09, 9.128476e-09, 9.118374e-09, 9.09953e-09, 9.118805e-09, 
    9.117238e-09, 9.135682e-09, 9.129755e-09, 9.174038e-09, 9.150251e-09, 
    9.217825e-09, 9.242485e-09, 9.312123e-09, 9.354813e-09, 9.398266e-09, 
    9.417451e-09, 9.423291e-09, 9.425731e-09 ;

 NFIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NFIX_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 OCDEP =
  3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14 ;

 O_SCALAR =
  0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 PARVEGLN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PBOT =
  102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8 ;

 PCH4 =
  0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993 ;

 PCO2 =
  29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676 ;

 PCT_LANDUNIT =
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PCT_NAT_PFT =
  13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892,
  55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_CTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_NTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PLANT_NDEMAND =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 POTENTIAL_IMMOB =
  4.490659e-14, 4.502776e-14, 4.500422e-14, 4.510187e-14, 4.504772e-14, 
    4.511163e-14, 4.493118e-14, 4.503255e-14, 4.496786e-14, 4.491753e-14, 
    4.529107e-14, 4.510622e-14, 4.548291e-14, 4.536523e-14, 4.566065e-14, 
    4.546458e-14, 4.570015e-14, 4.565504e-14, 4.579087e-14, 4.575198e-14, 
    4.592545e-14, 4.580882e-14, 4.601533e-14, 4.589763e-14, 4.591603e-14, 
    4.580496e-14, 4.514348e-14, 4.526806e-14, 4.513609e-14, 4.515386e-14, 
    4.51459e-14, 4.504883e-14, 4.499986e-14, 4.489735e-14, 4.491597e-14, 
    4.499127e-14, 4.516186e-14, 4.510401e-14, 4.524983e-14, 4.524654e-14, 
    4.540864e-14, 4.533558e-14, 4.560769e-14, 4.553044e-14, 4.57536e-14, 
    4.569751e-14, 4.575096e-14, 4.573476e-14, 4.575117e-14, 4.56689e-14, 
    4.570415e-14, 4.563174e-14, 4.534926e-14, 4.543234e-14, 4.518434e-14, 
    4.503489e-14, 4.493562e-14, 4.48651e-14, 4.487507e-14, 4.489407e-14, 
    4.499171e-14, 4.508348e-14, 4.515335e-14, 4.520005e-14, 4.524606e-14, 
    4.538511e-14, 4.545872e-14, 4.562329e-14, 4.559364e-14, 4.564389e-14, 
    4.569193e-14, 4.577248e-14, 4.575923e-14, 4.57947e-14, 4.564259e-14, 
    4.57437e-14, 4.557676e-14, 4.562242e-14, 4.525843e-14, 4.511962e-14, 
    4.506046e-14, 4.500874e-14, 4.488274e-14, 4.496976e-14, 4.493546e-14, 
    4.501708e-14, 4.506889e-14, 4.504327e-14, 4.520133e-14, 4.51399e-14, 
    4.546308e-14, 4.532399e-14, 4.568633e-14, 4.559973e-14, 4.570708e-14, 
    4.565232e-14, 4.574612e-14, 4.56617e-14, 4.580791e-14, 4.583971e-14, 
    4.581798e-14, 4.590147e-14, 4.565702e-14, 4.575095e-14, 4.504255e-14, 
    4.504672e-14, 4.50662e-14, 4.498056e-14, 4.497533e-14, 4.489683e-14, 
    4.496669e-14, 4.499642e-14, 4.50719e-14, 4.51165e-14, 4.515889e-14, 
    4.525204e-14, 4.535595e-14, 4.550115e-14, 4.560534e-14, 4.567514e-14, 
    4.563236e-14, 4.567013e-14, 4.56279e-14, 4.56081e-14, 4.582779e-14, 
    4.570447e-14, 4.588947e-14, 4.587924e-14, 4.579554e-14, 4.58804e-14, 
    4.504966e-14, 4.502562e-14, 4.494205e-14, 4.500745e-14, 4.488828e-14, 
    4.495499e-14, 4.499331e-14, 4.514116e-14, 4.517365e-14, 4.520372e-14, 
    4.526313e-14, 4.533932e-14, 4.547283e-14, 4.558886e-14, 4.569473e-14, 
    4.568698e-14, 4.56897e-14, 4.571333e-14, 4.565478e-14, 4.572294e-14, 
    4.573436e-14, 4.570447e-14, 4.587787e-14, 4.582837e-14, 4.587903e-14, 
    4.58468e-14, 4.503343e-14, 4.50739e-14, 4.505203e-14, 4.509313e-14, 
    4.506417e-14, 4.519288e-14, 4.523144e-14, 4.541174e-14, 4.533781e-14, 
    4.545548e-14, 4.534978e-14, 4.536851e-14, 4.545926e-14, 4.53555e-14, 
    4.558244e-14, 4.542859e-14, 4.571425e-14, 4.556073e-14, 4.572385e-14, 
    4.569427e-14, 4.574327e-14, 4.578711e-14, 4.584228e-14, 4.594395e-14, 
    4.592042e-14, 4.600542e-14, 4.51342e-14, 4.518662e-14, 4.518203e-14, 
    4.523689e-14, 4.527743e-14, 4.536528e-14, 4.550603e-14, 4.545313e-14, 
    4.555025e-14, 4.556973e-14, 4.542219e-14, 4.551277e-14, 4.522171e-14, 
    4.526876e-14, 4.524076e-14, 4.513832e-14, 4.546528e-14, 4.529759e-14, 
    4.560706e-14, 4.551639e-14, 4.578086e-14, 4.564937e-14, 4.590746e-14, 
    4.601754e-14, 4.612116e-14, 4.624199e-14, 4.521525e-14, 4.517964e-14, 
    4.524341e-14, 4.533154e-14, 4.541332e-14, 4.552192e-14, 4.553304e-14, 
    4.555336e-14, 4.560599e-14, 4.565023e-14, 4.555976e-14, 4.566132e-14, 
    4.527962e-14, 4.547984e-14, 4.516615e-14, 4.526067e-14, 4.532636e-14, 
    4.529757e-14, 4.544709e-14, 4.548229e-14, 4.562519e-14, 4.555137e-14, 
    4.599036e-14, 4.579634e-14, 4.633398e-14, 4.618399e-14, 4.516718e-14, 
    4.521514e-14, 4.538182e-14, 4.530255e-14, 4.552917e-14, 4.558485e-14, 
    4.563014e-14, 4.568796e-14, 4.569422e-14, 4.572846e-14, 4.567234e-14, 
    4.572626e-14, 4.552215e-14, 4.56134e-14, 4.536281e-14, 4.542384e-14, 
    4.539578e-14, 4.536497e-14, 4.546003e-14, 4.556118e-14, 4.556338e-14, 
    4.559576e-14, 4.568695e-14, 4.553009e-14, 4.60153e-14, 4.571581e-14, 
    4.52674e-14, 4.53596e-14, 4.537281e-14, 4.53371e-14, 4.557929e-14, 
    4.549159e-14, 4.572763e-14, 4.566389e-14, 4.576832e-14, 4.571644e-14, 
    4.57088e-14, 4.564213e-14, 4.560059e-14, 4.549561e-14, 4.541011e-14, 
    4.534228e-14, 4.535806e-14, 4.543255e-14, 4.556737e-14, 4.569476e-14, 
    4.566686e-14, 4.576039e-14, 4.551275e-14, 4.561662e-14, 4.557649e-14, 
    4.568115e-14, 4.545171e-14, 4.5647e-14, 4.540172e-14, 4.542326e-14, 
    4.548985e-14, 4.562364e-14, 4.565328e-14, 4.568485e-14, 4.566539e-14, 
    4.55708e-14, 4.555531e-14, 4.548824e-14, 4.54697e-14, 4.541857e-14, 
    4.537621e-14, 4.54149e-14, 4.545552e-14, 4.557085e-14, 4.567464e-14, 
    4.578773e-14, 4.581541e-14, 4.594725e-14, 4.583988e-14, 4.601695e-14, 
    4.586634e-14, 4.612697e-14, 4.565836e-14, 4.586199e-14, 4.549289e-14, 
    4.553273e-14, 4.560467e-14, 4.576966e-14, 4.568066e-14, 4.578475e-14, 
    4.555471e-14, 4.54351e-14, 4.540418e-14, 4.53464e-14, 4.540551e-14, 
    4.54007e-14, 4.545723e-14, 4.543907e-14, 4.557468e-14, 4.550186e-14, 
    4.570859e-14, 4.578394e-14, 4.59965e-14, 4.612657e-14, 4.625888e-14, 
    4.631722e-14, 4.633497e-14, 4.634239e-14 ;

 POT_F_DENIT =
  1.021991e-12, 1.024835e-12, 1.024281e-12, 1.026576e-12, 1.025302e-12, 
    1.026804e-12, 1.022565e-12, 1.024945e-12, 1.023425e-12, 1.022242e-12, 
    1.031023e-12, 1.026674e-12, 1.035533e-12, 1.032761e-12, 1.039718e-12, 
    1.035101e-12, 1.040648e-12, 1.039582e-12, 1.042783e-12, 1.041865e-12, 
    1.04596e-12, 1.043205e-12, 1.048079e-12, 1.045301e-12, 1.045735e-12, 
    1.043112e-12, 1.027552e-12, 1.030486e-12, 1.027377e-12, 1.027796e-12, 
    1.027607e-12, 1.025326e-12, 1.024178e-12, 1.021768e-12, 1.022205e-12, 
    1.023974e-12, 1.02798e-12, 1.026618e-12, 1.030044e-12, 1.029967e-12, 
    1.03378e-12, 1.032061e-12, 1.038466e-12, 1.036645e-12, 1.041903e-12, 
    1.04058e-12, 1.04184e-12, 1.041457e-12, 1.041844e-12, 1.039905e-12, 
    1.040735e-12, 1.039028e-12, 1.032389e-12, 1.034344e-12, 1.02851e-12, 
    1.025002e-12, 1.022667e-12, 1.021012e-12, 1.021245e-12, 1.021691e-12, 
    1.023983e-12, 1.026136e-12, 1.027777e-12, 1.028874e-12, 1.029954e-12, 
    1.03323e-12, 1.03496e-12, 1.038834e-12, 1.038133e-12, 1.039318e-12, 
    1.040448e-12, 1.042347e-12, 1.042034e-12, 1.04287e-12, 1.039283e-12, 
    1.041667e-12, 1.03773e-12, 1.038807e-12, 1.030258e-12, 1.026988e-12, 
    1.025601e-12, 1.024383e-12, 1.021424e-12, 1.023468e-12, 1.022662e-12, 
    1.024576e-12, 1.025793e-12, 1.02519e-12, 1.028903e-12, 1.027459e-12, 
    1.035062e-12, 1.031788e-12, 1.040317e-12, 1.038276e-12, 1.040804e-12, 
    1.039514e-12, 1.041725e-12, 1.039734e-12, 1.04318e-12, 1.043931e-12, 
    1.043417e-12, 1.045386e-12, 1.039621e-12, 1.041836e-12, 1.025176e-12, 
    1.025274e-12, 1.025731e-12, 1.023721e-12, 1.023597e-12, 1.021753e-12, 
    1.023392e-12, 1.024091e-12, 1.025861e-12, 1.026909e-12, 1.027904e-12, 
    1.030094e-12, 1.032539e-12, 1.035955e-12, 1.038408e-12, 1.040051e-12, 
    1.039042e-12, 1.039932e-12, 1.038937e-12, 1.038469e-12, 1.043648e-12, 
    1.040741e-12, 1.045101e-12, 1.04486e-12, 1.042886e-12, 1.044886e-12, 
    1.025342e-12, 1.024776e-12, 1.022815e-12, 1.024349e-12, 1.021551e-12, 
    1.023118e-12, 1.024018e-12, 1.027489e-12, 1.02825e-12, 1.028958e-12, 
    1.030354e-12, 1.032145e-12, 1.035287e-12, 1.038019e-12, 1.040512e-12, 
    1.040328e-12, 1.040392e-12, 1.040949e-12, 1.039569e-12, 1.041174e-12, 
    1.041444e-12, 1.040739e-12, 1.044826e-12, 1.043658e-12, 1.044853e-12, 
    1.044091e-12, 1.024959e-12, 1.025909e-12, 1.025395e-12, 1.026361e-12, 
    1.02568e-12, 1.028705e-12, 1.029612e-12, 1.033852e-12, 1.03211e-12, 
    1.03488e-12, 1.03239e-12, 1.032831e-12, 1.03497e-12, 1.032523e-12, 
    1.037868e-12, 1.034245e-12, 1.04097e-12, 1.037356e-12, 1.041195e-12, 
    1.040497e-12, 1.041651e-12, 1.042686e-12, 1.043985e-12, 1.046385e-12, 
    1.045828e-12, 1.047834e-12, 1.027325e-12, 1.028558e-12, 1.028448e-12, 
    1.029737e-12, 1.03069e-12, 1.032756e-12, 1.036068e-12, 1.034822e-12, 
    1.037107e-12, 1.037567e-12, 1.034092e-12, 1.036226e-12, 1.029377e-12, 
    1.030484e-12, 1.029823e-12, 1.027415e-12, 1.035106e-12, 1.03116e-12, 
    1.038442e-12, 1.036305e-12, 1.042537e-12, 1.039439e-12, 1.045522e-12, 
    1.048124e-12, 1.050566e-12, 1.053424e-12, 1.029229e-12, 1.028391e-12, 
    1.029889e-12, 1.031964e-12, 1.033885e-12, 1.036442e-12, 1.036702e-12, 
    1.037181e-12, 1.038419e-12, 1.039462e-12, 1.037331e-12, 1.039722e-12, 
    1.030742e-12, 1.035448e-12, 1.028068e-12, 1.030292e-12, 1.031834e-12, 
    1.031156e-12, 1.034672e-12, 1.035501e-12, 1.038867e-12, 1.037126e-12, 
    1.047481e-12, 1.042902e-12, 1.055595e-12, 1.052051e-12, 1.028098e-12, 
    1.029224e-12, 1.033145e-12, 1.031279e-12, 1.036611e-12, 1.037923e-12, 
    1.038988e-12, 1.040352e-12, 1.040497e-12, 1.041305e-12, 1.03998e-12, 
    1.041251e-12, 1.036442e-12, 1.038591e-12, 1.03269e-12, 1.034126e-12, 
    1.033465e-12, 1.032739e-12, 1.034975e-12, 1.037359e-12, 1.037408e-12, 
    1.038172e-12, 1.040328e-12, 1.036623e-12, 1.048072e-12, 1.041005e-12, 
    1.030452e-12, 1.032622e-12, 1.03293e-12, 1.03209e-12, 1.03779e-12, 
    1.035725e-12, 1.041285e-12, 1.039782e-12, 1.042243e-12, 1.04102e-12, 
    1.040839e-12, 1.039267e-12, 1.038288e-12, 1.035816e-12, 1.033802e-12, 
    1.032205e-12, 1.032576e-12, 1.03433e-12, 1.037504e-12, 1.040505e-12, 
    1.039847e-12, 1.042049e-12, 1.036214e-12, 1.038662e-12, 1.037715e-12, 
    1.04018e-12, 1.034787e-12, 1.039393e-12, 1.033609e-12, 1.034115e-12, 
    1.035682e-12, 1.038836e-12, 1.039531e-12, 1.040276e-12, 1.039815e-12, 
    1.037588e-12, 1.037221e-12, 1.035641e-12, 1.035204e-12, 1.034e-12, 
    1.033002e-12, 1.033913e-12, 1.034869e-12, 1.037584e-12, 1.04003e-12, 
    1.042694e-12, 1.043346e-12, 1.046461e-12, 1.043926e-12, 1.048109e-12, 
    1.044555e-12, 1.050704e-12, 1.039656e-12, 1.044458e-12, 1.035754e-12, 
    1.036691e-12, 1.038388e-12, 1.042276e-12, 1.040175e-12, 1.042631e-12, 
    1.037207e-12, 1.034392e-12, 1.033661e-12, 1.032302e-12, 1.033691e-12, 
    1.033578e-12, 1.034908e-12, 1.03448e-12, 1.037673e-12, 1.035957e-12, 
    1.040828e-12, 1.042605e-12, 1.047619e-12, 1.050691e-12, 1.053815e-12, 
    1.055193e-12, 1.055613e-12, 1.055787e-12 ;

 POT_F_NIT =
  4.014551e-11, 4.049193e-11, 4.042445e-11, 4.070474e-11, 4.054912e-11, 
    4.073283e-11, 4.021559e-11, 4.050569e-11, 4.032037e-11, 4.017659e-11, 
    4.125151e-11, 4.071723e-11, 4.181026e-11, 4.146671e-11, 4.233246e-11, 
    4.17567e-11, 4.244905e-11, 4.231578e-11, 4.27175e-11, 4.260221e-11, 
    4.31182e-11, 4.277076e-11, 4.338693e-11, 4.303508e-11, 4.309002e-11, 
    4.27593e-11, 4.082448e-11, 4.118484e-11, 4.080318e-11, 4.085445e-11, 
    4.083144e-11, 4.055232e-11, 4.041205e-11, 4.011905e-11, 4.017215e-11, 
    4.038738e-11, 4.087749e-11, 4.071076e-11, 4.113158e-11, 4.112206e-11, 
    4.159313e-11, 4.138039e-11, 4.21763e-11, 4.194928e-11, 4.260701e-11, 
    4.24411e-11, 4.25992e-11, 4.255122e-11, 4.259982e-11, 4.235663e-11, 
    4.246073e-11, 4.224705e-11, 4.142024e-11, 4.166238e-11, 4.094233e-11, 
    4.05125e-11, 4.022828e-11, 4.002723e-11, 4.005561e-11, 4.010977e-11, 
    4.038864e-11, 4.065173e-11, 4.085283e-11, 4.098763e-11, 4.112067e-11, 
    4.152479e-11, 4.173948e-11, 4.222228e-11, 4.213492e-11, 4.228295e-11, 
    4.24246e-11, 4.266299e-11, 4.26237e-11, 4.272889e-11, 4.227901e-11, 
    4.257773e-11, 4.208518e-11, 4.22196e-11, 4.115696e-11, 4.075572e-11, 
    4.058582e-11, 4.043738e-11, 4.007744e-11, 4.032583e-11, 4.022781e-11, 
    4.046117e-11, 4.060982e-11, 4.053626e-11, 4.099131e-11, 4.081408e-11, 
    4.175221e-11, 4.134678e-11, 4.240807e-11, 4.215283e-11, 4.246935e-11, 
    4.230769e-11, 4.258488e-11, 4.233536e-11, 4.276807e-11, 4.28626e-11, 
    4.279798e-11, 4.304643e-11, 4.232152e-11, 4.259916e-11, 4.053422e-11, 
    4.054622e-11, 4.06021e-11, 4.035672e-11, 4.034173e-11, 4.011757e-11, 
    4.031699e-11, 4.040206e-11, 4.061843e-11, 4.07467e-11, 4.086882e-11, 
    4.113801e-11, 4.143972e-11, 4.186352e-11, 4.216935e-11, 4.2375e-11, 
    4.224883e-11, 4.236021e-11, 4.22357e-11, 4.217741e-11, 4.282716e-11, 
    4.246168e-11, 4.301064e-11, 4.298017e-11, 4.273137e-11, 4.298359e-11, 
    4.055463e-11, 4.048563e-11, 4.024659e-11, 4.043359e-11, 4.009319e-11, 
    4.028355e-11, 4.039321e-11, 4.081778e-11, 4.091136e-11, 4.099825e-11, 
    4.117012e-11, 4.139123e-11, 4.178061e-11, 4.212092e-11, 4.243283e-11, 
    4.240993e-11, 4.241799e-11, 4.248782e-11, 4.231495e-11, 4.251622e-11, 
    4.255005e-11, 4.246162e-11, 4.297608e-11, 4.282877e-11, 4.297951e-11, 
    4.288355e-11, 4.050804e-11, 4.062419e-11, 4.05614e-11, 4.06795e-11, 
    4.059628e-11, 4.096701e-11, 4.10785e-11, 4.160226e-11, 4.138687e-11, 
    4.172991e-11, 4.142164e-11, 4.147618e-11, 4.174113e-11, 4.143826e-11, 
    4.210211e-11, 4.165145e-11, 4.249053e-11, 4.203836e-11, 4.251894e-11, 
    4.243145e-11, 4.257633e-11, 4.270632e-11, 4.287013e-11, 4.317326e-11, 
    4.310296e-11, 4.33571e-11, 4.079765e-11, 4.094889e-11, 4.093556e-11, 
    4.109411e-11, 4.121157e-11, 4.146675e-11, 4.187774e-11, 4.172293e-11, 
    4.200734e-11, 4.206455e-11, 4.163255e-11, 4.189752e-11, 4.105023e-11, 
    4.118651e-11, 4.110533e-11, 4.080952e-11, 4.175855e-11, 4.127009e-11, 
    4.217436e-11, 4.190802e-11, 4.268777e-11, 4.229906e-11, 4.306429e-11, 
    4.339361e-11, 4.370469e-11, 4.406973e-11, 4.103155e-11, 4.092864e-11, 
    4.111297e-11, 4.136873e-11, 4.160675e-11, 4.192429e-11, 4.195684e-11, 
    4.201649e-11, 4.217119e-11, 4.230151e-11, 4.203536e-11, 4.23342e-11, 
    4.121816e-11, 4.180109e-11, 4.088972e-11, 4.116307e-11, 4.135358e-11, 
    4.126994e-11, 4.170521e-11, 4.180813e-11, 4.222776e-11, 4.201057e-11, 
    4.33122e-11, 4.273379e-11, 4.434871e-11, 4.389429e-11, 4.089271e-11, 
    4.103117e-11, 4.151497e-11, 4.128441e-11, 4.194552e-11, 4.210909e-11, 
    4.224228e-11, 4.241289e-11, 4.243132e-11, 4.253259e-11, 4.236669e-11, 
    4.252602e-11, 4.192493e-11, 4.219299e-11, 4.145947e-11, 4.163739e-11, 
    4.155548e-11, 4.146574e-11, 4.174302e-11, 4.20395e-11, 4.204583e-11, 
    4.214112e-11, 4.24103e-11, 4.194813e-11, 4.338716e-11, 4.24955e-11, 
    4.118243e-11, 4.145034e-11, 4.148866e-11, 4.138473e-11, 4.209266e-11, 
    4.183543e-11, 4.253012e-11, 4.234178e-11, 4.265058e-11, 4.249698e-11, 
    4.24744e-11, 4.22776e-11, 4.215531e-11, 4.184718e-11, 4.159732e-11, 
    4.139974e-11, 4.144563e-11, 4.166282e-11, 4.205765e-11, 4.243294e-11, 
    4.235058e-11, 4.262701e-11, 4.189732e-11, 4.22025e-11, 4.208441e-11, 
    4.239267e-11, 4.171881e-11, 4.22924e-11, 4.157285e-11, 4.163567e-11, 
    4.183032e-11, 4.222332e-11, 4.231049e-11, 4.240371e-11, 4.234616e-11, 
    4.206773e-11, 4.202219e-11, 4.182556e-11, 4.177135e-11, 4.162195e-11, 
    4.149846e-11, 4.161127e-11, 4.172991e-11, 4.206781e-11, 4.237352e-11, 
    4.270813e-11, 4.279021e-11, 4.318331e-11, 4.286318e-11, 4.339213e-11, 
    4.294223e-11, 4.372255e-11, 4.232573e-11, 4.29291e-11, 4.183919e-11, 
    4.19559e-11, 4.216745e-11, 4.26547e-11, 4.239127e-11, 4.269943e-11, 
    4.20204e-11, 4.167034e-11, 4.157999e-11, 4.141174e-11, 4.158383e-11, 
    4.156982e-11, 4.173482e-11, 4.168175e-11, 4.207904e-11, 4.186539e-11, 
    4.247378e-11, 4.269694e-11, 4.333038e-11, 4.372109e-11, 4.412066e-11, 
    4.429766e-11, 4.435161e-11, 4.437416e-11 ;

 PROD100C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHADE_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Q2M =
  0.001208388, 0.001208317, 0.001208331, 0.001208274, 0.001208305, 
    0.001208268, 0.001208373, 0.001208315, 0.001208352, 0.001208381, 
    0.001208165, 0.001208271, 0.00120805, 0.001208118, 0.001207944, 
    0.001208062, 0.00120792, 0.001207946, 0.001207865, 0.001207888, 
    0.001207788, 0.001207855, 0.001207735, 0.001207804, 0.001207793, 
    0.001207857, 0.001208249, 0.001208179, 0.001208253, 0.001208243, 
    0.001208247, 0.001208305, 0.001208335, 0.001208393, 0.001208382, 
    0.001208339, 0.001208238, 0.001208272, 0.001208185, 0.001208187, 
    0.001208093, 0.001208135, 0.001207974, 0.00120802, 0.001207887, 
    0.001207921, 0.001207889, 0.001207899, 0.001207889, 0.001207938, 
    0.001207917, 0.001207959, 0.001208128, 0.001208079, 0.001208225, 
    0.001208315, 0.001208371, 0.001208412, 0.001208406, 0.001208396, 
    0.001208339, 0.001208284, 0.001208242, 0.001208215, 0.001208188, 
    0.001208109, 0.001208064, 0.001207965, 0.001207982, 0.001207953, 
    0.001207924, 0.001207877, 0.001207884, 0.001207864, 0.001207953, 
    0.001207894, 0.001207993, 0.001207965, 0.001208185, 0.001208262, 
    0.001208299, 0.001208328, 0.001208402, 0.001208351, 0.001208371, 
    0.001208323, 0.001208292, 0.001208307, 0.001208214, 0.00120825, 
    0.001208062, 0.001208143, 0.001207927, 0.001207978, 0.001207915, 
    0.001207947, 0.001207892, 0.001207942, 0.001207856, 0.001207838, 
    0.00120785, 0.001207801, 0.001207944, 0.00120789, 0.001208308, 
    0.001208305, 0.001208294, 0.001208345, 0.001208348, 0.001208394, 
    0.001208353, 0.001208335, 0.00120829, 0.001208264, 0.001208239, 
    0.001208185, 0.001208124, 0.001208039, 0.001207975, 0.001207934, 
    0.001207959, 0.001207937, 0.001207961, 0.001207973, 0.001207845, 
    0.001207917, 0.001207808, 0.001207814, 0.001207863, 0.001207813, 
    0.001208304, 0.001208317, 0.001208367, 0.001208328, 0.001208398, 
    0.00120836, 0.001208338, 0.001208251, 0.001208231, 0.001208213, 
    0.001208178, 0.001208133, 0.001208055, 0.001207985, 0.001207922, 
    0.001207927, 0.001207925, 0.001207911, 0.001207946, 0.001207906, 
    0.001207899, 0.001207917, 0.001207814, 0.001207843, 0.001207814, 
    0.001207832, 0.001208313, 0.001208289, 0.001208302, 0.001208278, 
    0.001208295, 0.00120822, 0.001208198, 0.001208092, 0.001208134, 
    0.001208066, 0.001208127, 0.001208116, 0.001208065, 0.001208123, 
    0.00120799, 0.001208083, 0.001207911, 0.001208005, 0.001207905, 
    0.001207922, 0.001207893, 0.001207868, 0.001207835, 0.001207776, 
    0.00120779, 0.00120774, 0.001208254, 0.001208224, 0.001208225, 
    0.001208193, 0.00120817, 0.001208118, 0.001208035, 0.001208066, 
    0.001208009, 0.001207998, 0.001208084, 0.001208032, 0.001208203, 
    0.001208176, 0.001208191, 0.001208252, 0.00120806, 0.001208159, 
    0.001207974, 0.001208029, 0.001207872, 0.00120795, 0.001207797, 
    0.001207735, 0.001207671, 0.001207602, 0.001208206, 0.001208227, 
    0.001208189, 0.001208139, 0.00120809, 0.001208026, 0.001208019, 
    0.001208007, 0.001207974, 0.001207948, 0.001208004, 0.001207942, 
    0.001208172, 0.001208051, 0.001208235, 0.001208181, 0.001208142, 
    0.001208158, 0.001208069, 0.001208049, 0.001207964, 0.001208008, 
    0.001207751, 0.001207864, 0.001207547, 0.001207636, 0.001208234, 
    0.001208206, 0.001208109, 0.001208155, 0.001208021, 0.001207987, 
    0.00120796, 0.001207927, 0.001207922, 0.001207903, 0.001207935, 
    0.001207904, 0.001208026, 0.00120797, 0.001208119, 0.001208084, 
    0.0012081, 0.001208118, 0.001208062, 0.001208004, 0.001208001, 
    0.001207981, 0.001207932, 0.001208021, 0.001207739, 0.001207914, 
    0.001208175, 0.001208123, 0.001208114, 0.001208134, 0.001207992, 
    0.001208044, 0.001207903, 0.00120794, 0.001207879, 0.001207909, 
    0.001207914, 0.001207953, 0.001207978, 0.001208042, 0.001208092, 
    0.001208131, 0.001208122, 0.001208079, 0.001208, 0.001207923, 
    0.001207939, 0.001207883, 0.001208031, 0.001207969, 0.001207994, 
    0.00120793, 0.001208067, 0.001207955, 0.001208096, 0.001208083, 
    0.001208045, 0.001207966, 0.001207946, 0.001207929, 0.001207939, 
    0.001207998, 0.001208006, 0.001208045, 0.001208057, 0.001208086, 
    0.001208111, 0.001208089, 0.001208065, 0.001207997, 0.001207935, 
    0.001207868, 0.001207851, 0.001207777, 0.001207839, 0.001207738, 
    0.001207827, 0.001207672, 0.001207946, 0.001207827, 0.001208042, 
    0.001208019, 0.001207976, 0.00120788, 0.001207931, 0.001207871, 
    0.001208007, 0.001208078, 0.001208095, 0.001208129, 0.001208094, 
    0.001208097, 0.001208063, 0.001208074, 0.001207995, 0.001208037, 
    0.001207914, 0.001207871, 0.001207746, 0.00120767, 0.00120759, 
    0.001207556, 0.001207546, 0.001207541 ;

 QBOT =
  0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224 ;

 QCHARGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_PERCH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_XS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRIP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLOOD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_ICE_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_LIQ_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINFL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QIRRIG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRGWL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QSNOMELT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSOIL =
  3.025561e-06, 3.032672e-06, 3.031294e-06, 3.037005e-06, 3.033852e-06, 
    3.037576e-06, 3.027012e-06, 3.032946e-06, 3.029163e-06, 3.026214e-06, 
    3.048023e-06, 3.037261e-06, 3.059291e-06, 3.052411e-06, 3.070438e-06, 
    3.058208e-06, 3.07277e-06, 3.070126e-06, 3.078138e-06, 3.075844e-06, 
    3.086055e-06, 3.079198e-06, 3.091387e-06, 3.084428e-06, 3.085508e-06, 
    3.078968e-06, 3.039446e-06, 3.046677e-06, 3.039014e-06, 3.040045e-06, 
    3.039587e-06, 3.03391e-06, 3.031019e-06, 3.025033e-06, 3.026123e-06, 
    3.030528e-06, 3.04051e-06, 3.037144e-06, 3.04567e-06, 3.045478e-06, 
    3.054955e-06, 3.05068e-06, 3.06734e-06, 3.062104e-06, 3.07594e-06, 
    3.07263e-06, 3.075781e-06, 3.074828e-06, 3.075793e-06, 3.070941e-06, 
    3.073018e-06, 3.068757e-06, 3.051477e-06, 3.056339e-06, 3.041829e-06, 
    3.033064e-06, 3.027269e-06, 3.023141e-06, 3.023724e-06, 3.024832e-06, 
    3.030553e-06, 3.035946e-06, 3.040029e-06, 3.042758e-06, 3.04545e-06, 
    3.053542e-06, 3.057873e-06, 3.068247e-06, 3.066517e-06, 3.069462e-06, 
    3.072302e-06, 3.077048e-06, 3.076269e-06, 3.078357e-06, 3.069397e-06, 
    3.075344e-06, 3.064827e-06, 3.068209e-06, 3.046111e-06, 3.038055e-06, 
    3.03457e-06, 3.031557e-06, 3.024171e-06, 3.029267e-06, 3.027256e-06, 
    3.032056e-06, 3.035093e-06, 3.033596e-06, 3.042833e-06, 3.03924e-06, 
    3.05813e-06, 3.049993e-06, 3.07197e-06, 3.066874e-06, 3.073196e-06, 
    3.069972e-06, 3.07549e-06, 3.070524e-06, 3.07914e-06, 3.081009e-06, 
    3.07973e-06, 3.084667e-06, 3.070247e-06, 3.075774e-06, 3.03355e-06, 
    3.033794e-06, 3.034939e-06, 3.029899e-06, 3.029595e-06, 3.024999e-06, 
    3.029095e-06, 3.030834e-06, 3.035274e-06, 3.037872e-06, 3.040348e-06, 
    3.045794e-06, 3.05186e-06, 3.060371e-06, 3.067203e-06, 3.071316e-06, 
    3.068798e-06, 3.07102e-06, 3.068534e-06, 3.067372e-06, 3.080304e-06, 
    3.073033e-06, 3.083957e-06, 3.083355e-06, 3.078404e-06, 3.083423e-06, 
    3.033967e-06, 3.032559e-06, 3.027648e-06, 3.031491e-06, 3.0245e-06, 
    3.028403e-06, 3.030643e-06, 3.0393e-06, 3.041214e-06, 3.042967e-06, 
    3.046445e-06, 3.050898e-06, 3.058712e-06, 3.066228e-06, 3.07247e-06, 
    3.072014e-06, 3.072174e-06, 3.073562e-06, 3.070114e-06, 3.074128e-06, 
    3.074796e-06, 3.073041e-06, 3.083274e-06, 3.08035e-06, 3.083342e-06, 
    3.08144e-06, 3.033019e-06, 3.035386e-06, 3.034108e-06, 3.036505e-06, 
    3.034813e-06, 3.042318e-06, 3.044569e-06, 3.05512e-06, 3.050807e-06, 
    3.057692e-06, 3.051512e-06, 3.052603e-06, 3.057886e-06, 3.05185e-06, 
    3.065837e-06, 3.0561e-06, 3.073616e-06, 3.063845e-06, 3.074183e-06, 
    3.072443e-06, 3.075331e-06, 3.077911e-06, 3.08117e-06, 3.087167e-06, 
    3.085781e-06, 3.09081e-06, 3.038908e-06, 3.041961e-06, 3.041705e-06, 
    3.04491e-06, 3.047277e-06, 3.052422e-06, 3.060664e-06, 3.057568e-06, 
    3.063268e-06, 3.064407e-06, 3.055757e-06, 3.061054e-06, 3.044014e-06, 
    3.046753e-06, 3.045133e-06, 3.039141e-06, 3.058263e-06, 3.04844e-06, 
    3.067302e-06, 3.061275e-06, 3.077541e-06, 3.06978e-06, 3.085015e-06, 
    3.091501e-06, 3.097673e-06, 3.104818e-06, 3.043642e-06, 3.041565e-06, 
    3.045295e-06, 3.050428e-06, 3.05523e-06, 3.061597e-06, 3.062256e-06, 
    3.063446e-06, 3.067247e-06, 3.069848e-06, 3.063809e-06, 3.070502e-06, 
    3.047361e-06, 3.059122e-06, 3.040768e-06, 3.046277e-06, 3.050131e-06, 
    3.048454e-06, 3.057218e-06, 3.05928e-06, 3.068362e-06, 3.063334e-06, 
    3.089888e-06, 3.078437e-06, 3.110307e-06, 3.10138e-06, 3.040837e-06, 
    3.043641e-06, 3.053377e-06, 3.048747e-06, 3.062029e-06, 3.065997e-06, 
    3.068668e-06, 3.072061e-06, 3.072438e-06, 3.074451e-06, 3.071151e-06, 
    3.074326e-06, 3.061611e-06, 3.067679e-06, 3.05228e-06, 3.055847e-06, 
    3.054211e-06, 3.052406e-06, 3.057975e-06, 3.063889e-06, 3.064037e-06, 
    3.066633e-06, 3.071938e-06, 3.062084e-06, 3.091327e-06, 3.073648e-06, 
    3.046697e-06, 3.052066e-06, 3.052859e-06, 3.050774e-06, 3.064968e-06, 
    3.05982e-06, 3.074405e-06, 3.070653e-06, 3.076808e-06, 3.073747e-06, 
    3.073296e-06, 3.069372e-06, 3.066924e-06, 3.060052e-06, 3.05504e-06, 
    3.051079e-06, 3.052002e-06, 3.056354e-06, 3.064256e-06, 3.072462e-06, 
    3.070814e-06, 3.07634e-06, 3.061065e-06, 3.06786e-06, 3.064795e-06, 
    3.071666e-06, 3.057481e-06, 3.069596e-06, 3.054559e-06, 3.05582e-06, 
    3.059718e-06, 3.068259e-06, 3.070028e-06, 3.071879e-06, 3.070741e-06, 
    3.064461e-06, 3.063558e-06, 3.059628e-06, 3.058533e-06, 3.055547e-06, 
    3.053065e-06, 3.055327e-06, 3.057699e-06, 3.064472e-06, 3.071276e-06, 
    3.077944e-06, 3.079585e-06, 3.08733e-06, 3.080995e-06, 3.091421e-06, 
    3.08251e-06, 3.097963e-06, 3.07029e-06, 3.082293e-06, 3.059902e-06, 
    3.06224e-06, 3.067148e-06, 3.07686e-06, 3.071637e-06, 3.077756e-06, 
    3.063524e-06, 3.056494e-06, 3.054702e-06, 3.051316e-06, 3.054779e-06, 
    3.054499e-06, 3.057812e-06, 3.056749e-06, 3.064698e-06, 3.060428e-06, 
    3.073278e-06, 3.077713e-06, 3.090275e-06, 3.097972e-06, 3.105849e-06, 
    3.109318e-06, 3.110376e-06, 3.110817e-06 ;

 QVEGE =
  -6.482299e-07, -6.477903e-07, -6.478738e-07, -6.475231e-07, -6.477144e-07, 
    -6.47487e-07, -6.481369e-07, -6.477764e-07, -6.480043e-07, -6.481849e-07, 
    -6.468516e-07, -6.475064e-07, -6.461357e-07, -6.465585e-07, 
    -6.454831e-07, -6.46207e-07, -6.453341e-07, -6.454948e-07, -6.449874e-07, 
    -6.451326e-07, -6.444996e-07, -6.449203e-07, -6.441542e-07, 
    -6.445953e-07, -6.4453e-07, -6.449357e-07, -6.473659e-07, -6.469356e-07, 
    -6.473934e-07, -6.473317e-07, -6.473574e-07, -6.477136e-07, 
    -6.478986e-07, -6.482572e-07, -6.481905e-07, -6.479237e-07, 
    -6.473037e-07, -6.475086e-07, -6.469733e-07, -6.469852e-07, 
    -6.463992e-07, -6.466638e-07, -6.4567e-07, -6.4595e-07, -6.451263e-07, 
    -6.453362e-07, -6.451378e-07, -6.451968e-07, -6.45137e-07, -6.454441e-07, 
    -6.453132e-07, -6.455799e-07, -6.466161e-07, -6.463148e-07, 
    -6.472188e-07, -6.477767e-07, -6.481228e-07, -6.483744e-07, 
    -6.483389e-07, -6.48273e-07, -6.479223e-07, -6.475834e-07, -6.473272e-07, 
    -6.471567e-07, -6.469871e-07, -6.465019e-07, -6.462242e-07, 
    -6.456173e-07, -6.457199e-07, -6.455401e-07, -6.453567e-07, 
    -6.450585e-07, -6.451065e-07, -6.449768e-07, -6.455391e-07, 
    -6.451687e-07, -6.457779e-07, -6.456143e-07, -6.469723e-07, 
    -6.474519e-07, -6.476816e-07, -6.478589e-07, -6.483122e-07, 
    -6.480011e-07, -6.481246e-07, -6.47824e-07, -6.476369e-07, -6.477282e-07, 
    -6.47152e-07, -6.473776e-07, -6.462078e-07, -6.467107e-07, -6.45378e-07, 
    -6.456982e-07, -6.453e-07, -6.455019e-07, -6.451582e-07, -6.454675e-07, 
    -6.449259e-07, -6.448111e-07, -6.448902e-07, -6.44575e-07, -6.454854e-07, 
    -6.451408e-07, -6.477322e-07, -6.477175e-07, -6.476454e-07, 
    -6.479626e-07, -6.479802e-07, -6.482605e-07, -6.480083e-07, 
    -6.479032e-07, -6.476236e-07, -6.474637e-07, -6.473092e-07, 
    -6.469683e-07, -6.465959e-07, -6.460643e-07, -6.456778e-07, 
    -6.454175e-07, -6.455751e-07, -6.454363e-07, -6.455927e-07, 
    -6.456646e-07, -6.448562e-07, -6.453138e-07, -6.446205e-07, 
    -6.446579e-07, -6.449749e-07, -6.446537e-07, -6.477067e-07, 
    -6.477922e-07, -6.480985e-07, -6.478588e-07, -6.482906e-07, 
    -6.480531e-07, -6.479185e-07, -6.473797e-07, -6.472534e-07, -6.47146e-07, 
    -6.469264e-07, -6.466504e-07, -6.46167e-07, -6.457416e-07, -6.453447e-07, 
    -6.453732e-07, -6.453635e-07, -6.452778e-07, -6.454942e-07, 
    -6.452419e-07, -6.452025e-07, -6.453102e-07, -6.446631e-07, 
    -6.448482e-07, -6.446588e-07, -6.447785e-07, -6.477636e-07, 
    -6.476182e-07, -6.476973e-07, -6.475502e-07, -6.476563e-07, 
    -6.471925e-07, -6.47053e-07, -6.463956e-07, -6.466576e-07, -6.462317e-07, 
    -6.46612e-07, -6.465465e-07, -6.462309e-07, -6.465895e-07, -6.457713e-07, 
    -6.463376e-07, -6.452744e-07, -6.458563e-07, -6.452384e-07, 
    -6.453465e-07, -6.451643e-07, -6.450043e-07, -6.447967e-07, 
    -6.444213e-07, -6.445071e-07, -6.441869e-07, -6.473981e-07, 
    -6.472115e-07, -6.472222e-07, -6.470223e-07, -6.468766e-07, 
    -6.465544e-07, -6.460427e-07, -6.462334e-07, -6.458766e-07, 
    -6.458068e-07, -6.463455e-07, -6.460207e-07, -6.470819e-07, -6.46916e-07, 
    -6.470102e-07, -6.473869e-07, -6.461976e-07, -6.468104e-07, 
    -6.456725e-07, -6.460033e-07, -6.45028e-07, -6.455218e-07, -6.445557e-07, 
    -6.441544e-07, -6.437471e-07, -6.433009e-07, -6.471031e-07, 
    -6.472308e-07, -6.469968e-07, -6.466864e-07, -6.463815e-07, 
    -6.459842e-07, -6.459402e-07, -6.458673e-07, -6.456728e-07, 
    -6.455101e-07, -6.458499e-07, -6.454686e-07, -6.468895e-07, 
    -6.461416e-07, -6.472844e-07, -6.469468e-07, -6.467021e-07, 
    -6.468034e-07, -6.462537e-07, -6.46126e-07, -6.456087e-07, -6.458723e-07, 
    -6.442589e-07, -6.449788e-07, -6.429394e-07, -6.435187e-07, 
    -6.472767e-07, -6.471008e-07, -6.465002e-07, -6.467844e-07, 
    -6.459545e-07, -6.457537e-07, -6.455833e-07, -6.453745e-07, 
    -6.453477e-07, -6.452228e-07, -6.454279e-07, -6.452287e-07, 
    -6.459834e-07, -6.456473e-07, -6.465618e-07, -6.463429e-07, 
    -6.464417e-07, -6.465542e-07, -6.462072e-07, -6.45846e-07, -6.458288e-07, 
    -6.457163e-07, -6.454092e-07, -6.459509e-07, -6.44183e-07, -6.452976e-07, 
    -6.469098e-07, -6.465863e-07, -6.465286e-07, -6.46656e-07, -6.457723e-07, 
    -6.460946e-07, -6.452245e-07, -6.454593e-07, -6.450718e-07, 
    -6.452654e-07, -6.452943e-07, -6.4554e-07, -6.456951e-07, -6.460817e-07, 
    -6.46394e-07, -6.466364e-07, -6.465793e-07, -6.463127e-07, -6.458217e-07, 
    -6.453494e-07, -6.454549e-07, -6.451012e-07, -6.460153e-07, 
    -6.456395e-07, -6.457868e-07, -6.45397e-07, -6.462406e-07, -6.455517e-07, 
    -6.464198e-07, -6.463418e-07, -6.461009e-07, -6.456201e-07, 
    -6.454987e-07, -6.45386e-07, -6.454536e-07, -6.458074e-07, -6.458613e-07, 
    -6.461045e-07, -6.461761e-07, -6.463581e-07, -6.46513e-07, -6.463738e-07, 
    -6.462295e-07, -6.458033e-07, -6.454244e-07, -6.450035e-07, 
    -6.448964e-07, -6.444247e-07, -6.44822e-07, -6.441787e-07, -6.447458e-07, 
    -6.437515e-07, -6.454976e-07, -6.447431e-07, -6.460868e-07, 
    -6.459408e-07, -6.45688e-07, -6.450796e-07, -6.453987e-07, -6.450207e-07, 
    -6.458627e-07, -6.463082e-07, -6.464115e-07, -6.466234e-07, 
    -6.464067e-07, -6.46424e-07, -6.462168e-07, -6.462828e-07, -6.45789e-07, 
    -6.460543e-07, -6.452976e-07, -6.450214e-07, -6.44224e-07, -6.437371e-07, 
    -6.432228e-07, -6.43e-07, -6.429311e-07, -6.429029e-07 ;

 QVEGT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RETRANSN =
  4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07 ;

 RETRANSN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RH2M =
  84.71109, 84.71064, 84.71072, 84.71038, 84.71057, 84.71035, 84.71099, 
    84.71062, 84.71086, 84.71104, 84.70976, 84.71037, 84.70921, 84.70954, 
    84.70829, 84.70926, 84.70818, 84.7083, 84.70795, 84.70805, 84.7076, 
    84.7079, 84.70738, 84.70767, 84.70763, 84.70791, 84.71024, 84.70984, 
    84.71027, 84.71021, 84.71023, 84.71056, 84.71075, 84.71112, 84.71105, 
    84.71078, 84.71018, 84.71037, 84.70988, 84.70989, 84.70941, 84.70963, 
    84.70843, 84.70908, 84.70804, 84.70819, 84.70805, 84.70809, 84.70805, 
    84.70827, 84.70817, 84.70836, 84.70959, 84.70935, 84.7101, 84.71062, 
    84.71098, 84.71124, 84.7112, 84.71114, 84.71078, 84.71044, 84.71021, 
    84.71004, 84.70989, 84.70949, 84.70927, 84.70838, 84.70847, 84.70833, 
    84.7082, 84.70799, 84.70802, 84.70793, 84.70834, 84.70807, 84.70895, 
    84.70839, 84.70987, 84.71032, 84.71053, 84.71071, 84.71117, 84.71085, 
    84.71098, 84.71068, 84.71049, 84.71059, 84.71004, 84.71025, 84.70927, 
    84.70966, 84.70821, 84.70845, 84.70816, 84.70831, 84.70806, 84.70828, 
    84.7079, 84.70782, 84.70788, 84.70766, 84.7083, 84.70805, 84.71059, 
    84.71057, 84.7105, 84.71082, 84.71083, 84.71112, 84.71086, 84.71075, 
    84.71048, 84.71033, 84.71019, 84.70988, 84.70957, 84.70916, 84.70844, 
    84.70824, 84.70836, 84.70826, 84.70837, 84.70843, 84.70785, 84.70817, 
    84.7077, 84.70772, 84.70793, 84.70772, 84.71056, 84.71065, 84.71095, 
    84.71072, 84.71115, 84.71091, 84.71077, 84.71025, 84.71014, 84.71004, 
    84.70984, 84.70962, 84.70924, 84.70847, 84.70819, 84.70821, 84.70821, 
    84.70815, 84.7083, 84.70812, 84.70809, 84.70817, 84.70773, 84.70785, 
    84.70772, 84.7078, 84.71062, 84.71048, 84.71056, 84.71041, 84.71051, 
    84.71008, 84.70995, 84.70941, 84.70962, 84.70928, 84.70959, 84.70953, 
    84.70927, 84.70956, 84.7085, 84.70937, 84.70815, 84.709, 84.70811, 
    84.7082, 84.70807, 84.70795, 84.70781, 84.70756, 84.70762, 84.70741, 
    84.71027, 84.7101, 84.71011, 84.70992, 84.7098, 84.70954, 84.70914, 
    84.70929, 84.70902, 84.70897, 84.70937, 84.70912, 84.70998, 84.70983, 
    84.70992, 84.71026, 84.70926, 84.70974, 84.70843, 84.70911, 84.70797, 
    84.70832, 84.70765, 84.70738, 84.70713, 84.70686, 84.71, 84.71011, 
    84.7099, 84.70964, 84.7094, 84.7091, 84.70907, 84.70901, 84.70843, 
    84.70831, 84.709, 84.70828, 84.7098, 84.70921, 84.71017, 84.70985, 
    84.70966, 84.70974, 84.7093, 84.70921, 84.70838, 84.70902, 84.70745, 
    84.70793, 84.70664, 84.70699, 84.71016, 84.71, 84.7095, 84.70972, 
    84.70908, 84.70849, 84.70837, 84.70821, 84.7082, 84.70811, 84.70825, 
    84.70811, 84.7091, 84.70841, 84.70955, 84.70937, 84.70945, 84.70954, 
    84.70927, 84.70899, 84.70898, 84.70846, 84.70822, 84.70908, 84.70739, 
    84.70815, 84.70983, 84.70956, 84.70952, 84.70962, 84.70895, 84.70918, 
    84.70811, 84.70827, 84.708, 84.70814, 84.70816, 84.70834, 84.70844, 
    84.70918, 84.70941, 84.7096, 84.70956, 84.70935, 84.70898, 84.7082, 
    84.70827, 84.70802, 84.70912, 84.7084, 84.70895, 84.70823, 84.70929, 
    84.70833, 84.70943, 84.70937, 84.70919, 84.70839, 84.70831, 84.70822, 
    84.70827, 84.70897, 84.70901, 84.70919, 84.70924, 84.70939, 84.7095, 
    84.7094, 84.70928, 84.70897, 84.70825, 84.70795, 84.70788, 84.70756, 
    84.70782, 84.70739, 84.70776, 84.70712, 84.7083, 84.70776, 84.70918, 
    84.70907, 84.70844, 84.708, 84.70823, 84.70796, 84.70901, 84.70934, 
    84.70943, 84.70959, 84.70942, 84.70943, 84.70927, 84.70933, 84.70895, 
    84.70915, 84.70816, 84.70796, 84.70743, 84.70712, 84.70681, 84.70668, 
    84.70664, 84.70663 ;

 RH2M_R =
  84.71109, 84.71064, 84.71072, 84.71038, 84.71057, 84.71035, 84.71099, 
    84.71062, 84.71086, 84.71104, 84.70976, 84.71037, 84.70921, 84.70954, 
    84.70829, 84.70926, 84.70818, 84.7083, 84.70795, 84.70805, 84.7076, 
    84.7079, 84.70738, 84.70767, 84.70763, 84.70791, 84.71024, 84.70984, 
    84.71027, 84.71021, 84.71023, 84.71056, 84.71075, 84.71112, 84.71105, 
    84.71078, 84.71018, 84.71037, 84.70988, 84.70989, 84.70941, 84.70963, 
    84.70843, 84.70908, 84.70804, 84.70819, 84.70805, 84.70809, 84.70805, 
    84.70827, 84.70817, 84.70836, 84.70959, 84.70935, 84.7101, 84.71062, 
    84.71098, 84.71124, 84.7112, 84.71114, 84.71078, 84.71044, 84.71021, 
    84.71004, 84.70989, 84.70949, 84.70927, 84.70838, 84.70847, 84.70833, 
    84.7082, 84.70799, 84.70802, 84.70793, 84.70834, 84.70807, 84.70895, 
    84.70839, 84.70987, 84.71032, 84.71053, 84.71071, 84.71117, 84.71085, 
    84.71098, 84.71068, 84.71049, 84.71059, 84.71004, 84.71025, 84.70927, 
    84.70966, 84.70821, 84.70845, 84.70816, 84.70831, 84.70806, 84.70828, 
    84.7079, 84.70782, 84.70788, 84.70766, 84.7083, 84.70805, 84.71059, 
    84.71057, 84.7105, 84.71082, 84.71083, 84.71112, 84.71086, 84.71075, 
    84.71048, 84.71033, 84.71019, 84.70988, 84.70957, 84.70916, 84.70844, 
    84.70824, 84.70836, 84.70826, 84.70837, 84.70843, 84.70785, 84.70817, 
    84.7077, 84.70772, 84.70793, 84.70772, 84.71056, 84.71065, 84.71095, 
    84.71072, 84.71115, 84.71091, 84.71077, 84.71025, 84.71014, 84.71004, 
    84.70984, 84.70962, 84.70924, 84.70847, 84.70819, 84.70821, 84.70821, 
    84.70815, 84.7083, 84.70812, 84.70809, 84.70817, 84.70773, 84.70785, 
    84.70772, 84.7078, 84.71062, 84.71048, 84.71056, 84.71041, 84.71051, 
    84.71008, 84.70995, 84.70941, 84.70962, 84.70928, 84.70959, 84.70953, 
    84.70927, 84.70956, 84.7085, 84.70937, 84.70815, 84.709, 84.70811, 
    84.7082, 84.70807, 84.70795, 84.70781, 84.70756, 84.70762, 84.70741, 
    84.71027, 84.7101, 84.71011, 84.70992, 84.7098, 84.70954, 84.70914, 
    84.70929, 84.70902, 84.70897, 84.70937, 84.70912, 84.70998, 84.70983, 
    84.70992, 84.71026, 84.70926, 84.70974, 84.70843, 84.70911, 84.70797, 
    84.70832, 84.70765, 84.70738, 84.70713, 84.70686, 84.71, 84.71011, 
    84.7099, 84.70964, 84.7094, 84.7091, 84.70907, 84.70901, 84.70843, 
    84.70831, 84.709, 84.70828, 84.7098, 84.70921, 84.71017, 84.70985, 
    84.70966, 84.70974, 84.7093, 84.70921, 84.70838, 84.70902, 84.70745, 
    84.70793, 84.70664, 84.70699, 84.71016, 84.71, 84.7095, 84.70972, 
    84.70908, 84.70849, 84.70837, 84.70821, 84.7082, 84.70811, 84.70825, 
    84.70811, 84.7091, 84.70841, 84.70955, 84.70937, 84.70945, 84.70954, 
    84.70927, 84.70899, 84.70898, 84.70846, 84.70822, 84.70908, 84.70739, 
    84.70815, 84.70983, 84.70956, 84.70952, 84.70962, 84.70895, 84.70918, 
    84.70811, 84.70827, 84.708, 84.70814, 84.70816, 84.70834, 84.70844, 
    84.70918, 84.70941, 84.7096, 84.70956, 84.70935, 84.70898, 84.7082, 
    84.70827, 84.70802, 84.70912, 84.7084, 84.70895, 84.70823, 84.70929, 
    84.70833, 84.70943, 84.70937, 84.70919, 84.70839, 84.70831, 84.70822, 
    84.70827, 84.70897, 84.70901, 84.70919, 84.70924, 84.70939, 84.7095, 
    84.7094, 84.70928, 84.70897, 84.70825, 84.70795, 84.70788, 84.70756, 
    84.70782, 84.70739, 84.70776, 84.70712, 84.7083, 84.70776, 84.70918, 
    84.70907, 84.70844, 84.708, 84.70823, 84.70796, 84.70901, 84.70934, 
    84.70943, 84.70959, 84.70942, 84.70943, 84.70927, 84.70933, 84.70895, 
    84.70915, 84.70816, 84.70796, 84.70743, 84.70712, 84.70681, 84.70668, 
    84.70664, 84.70663 ;

 RH2M_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 RR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABG =
  0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 0.03212643, 
    0.03212643, 0.03212643 ;

 SABG_PEN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN =
  0.0004631664, 0.0004651067, 0.0004647294, 0.0004662944, 0.0004654261, 
    0.0004664508, 0.0004635594, 0.0004651835, 0.0004641466, 0.0004633405, 
    0.000469331, 0.0004663637, 0.0004724115, 0.0004705196, 0.0004752712, 
    0.0004721171, 0.000475907, 0.0004751798, 0.0004773675, 0.0004767407, 
    0.000479539, 0.0004776566, 0.000480989, 0.0004790893, 0.0004793865, 
    0.0004775943, 0.0004669611, 0.000468962, 0.0004668424, 0.0004671278, 
    0.0004669997, 0.0004654439, 0.00046466, 0.0004630174, 0.0004633155, 
    0.0004645218, 0.0004672557, 0.0004663274, 0.0004686661, 0.0004686132, 
    0.0004712165, 0.0004700428, 0.0004744177, 0.0004731742, 0.0004767668, 
    0.0004758633, 0.0004767243, 0.0004764631, 0.0004767276, 0.0004754026, 
    0.0004759702, 0.0004748042, 0.0004702633, 0.0004715983, 0.0004676162, 
    0.0004652217, 0.0004636305, 0.0004625015, 0.0004626609, 0.0004629653, 
    0.0004645287, 0.0004659984, 0.0004671183, 0.0004678674, 0.0004686055, 
    0.0004708402, 0.0004720222, 0.0004746691, 0.0004741912, 0.0004750005, 
    0.0004757734, 0.0004770711, 0.0004768574, 0.0004774292, 0.0004749787, 
    0.0004766074, 0.0004739186, 0.0004746541, 0.0004688075, 0.0004665781, 
    0.0004656311, 0.0004648014, 0.0004627836, 0.0004641771, 0.0004636278, 
    0.0004649343, 0.0004657645, 0.0004653538, 0.0004678879, 0.0004669027, 
    0.0004720922, 0.000469857, 0.0004756833, 0.0004742891, 0.0004760172, 
    0.0004751354, 0.0004766463, 0.0004752864, 0.0004776418, 0.0004781548, 
    0.0004778041, 0.0004791503, 0.0004752107, 0.0004767238, 0.0004653426, 
    0.0004654096, 0.0004657215, 0.0004643501, 0.0004642661, 0.000463009, 
    0.0004641273, 0.0004646037, 0.0004658125, 0.0004665275, 0.0004672071, 
    0.0004687015, 0.0004703704, 0.0004727036, 0.0004743795, 0.0004755027, 
    0.0004748139, 0.000475422, 0.0004747421, 0.0004744233, 0.0004779625, 
    0.0004759753, 0.0004789566, 0.0004787916, 0.0004774424, 0.00047881, 
    0.0004654565, 0.000465071, 0.000463733, 0.00046478, 0.0004628719, 
    0.0004639401, 0.0004645542, 0.0004669233, 0.0004674436, 0.0004679263, 
    0.0004688793, 0.0004701024, 0.000472248, 0.0004741145, 0.0004758181, 
    0.0004756932, 0.0004757371, 0.0004761177, 0.0004751749, 0.0004762723, 
    0.0004764565, 0.0004759748, 0.0004787693, 0.000477971, 0.0004787878, 
    0.0004782679, 0.0004651962, 0.0004658446, 0.0004654941, 0.0004661531, 
    0.0004656888, 0.000467753, 0.0004683718, 0.0004712668, 0.0004700784, 
    0.0004719694, 0.0004702703, 0.0004705714, 0.0004720312, 0.0004703619, 
    0.0004740116, 0.0004715375, 0.0004761324, 0.0004736624, 0.0004762871, 
    0.0004758103, 0.0004765994, 0.0004773063, 0.0004781952, 0.0004798358, 
    0.0004794557, 0.0004808276, 0.0004668112, 0.0004676523, 0.0004675781, 
    0.0004684581, 0.0004691089, 0.0004705194, 0.0004727816, 0.0004719308, 
    0.0004734923, 0.0004738058, 0.0004714332, 0.0004728901, 0.0004682145, 
    0.0004689701, 0.00046852, 0.0004668768, 0.0004721266, 0.0004694326, 
    0.0004744066, 0.0004729473, 0.0004772053, 0.000475088, 0.0004792466, 
    0.0004810246, 0.0004826968, 0.0004846518, 0.0004681111, 0.0004675395, 
    0.0004685626, 0.0004699783, 0.0004712913, 0.000473037, 0.0004732154, 
    0.0004735424, 0.0004743893, 0.0004751015, 0.0004736459, 0.0004752799, 
    0.0004691456, 0.0004723603, 0.0004673229, 0.0004688401, 0.0004698941, 
    0.0004694315, 0.0004718328, 0.0004723987, 0.0004746984, 0.0004735095, 
    0.0004805857, 0.0004774554, 0.0004861396, 0.0004837133, 0.0004673398, 
    0.0004681088, 0.0004707855, 0.0004695119, 0.0004731533, 0.0004740496, 
    0.0004747779, 0.0004757093, 0.0004758096, 0.0004763615, 0.0004754571, 
    0.0004763256, 0.0004730401, 0.0004745084, 0.0004704788, 0.0004714596, 
    0.0004710083, 0.0004705132, 0.0004720407, 0.0004736682, 0.0004737026, 
    0.0004742244, 0.0004756954, 0.000473167, 0.00048099, 0.0004761595, 
    0.0004689474, 0.0004704289, 0.0004706402, 0.0004700663, 0.0004739596, 
    0.000472549, 0.000476348, 0.0004753212, 0.0004770033, 0.0004761674, 
    0.0004760443, 0.0004749707, 0.0004743022, 0.0004726133, 0.0004712389, 
    0.0004701489, 0.0004704022, 0.0004715995, 0.0004737675, 0.0004758182, 
    0.000475369, 0.0004768747, 0.0004728882, 0.00047456, 0.0004739139, 
    0.0004755984, 0.000471908, 0.0004750524, 0.0004711042, 0.0004714503, 
    0.0004725209, 0.0004746745, 0.0004751504, 0.0004756591, 0.000475345, 
    0.0004738229, 0.0004735734, 0.0004724944, 0.0004721966, 0.0004713744, 
    0.0004706937, 0.0004713156, 0.0004719686, 0.000473823, 0.0004754941, 
    0.0004773157, 0.0004777613, 0.00047989, 0.0004781575, 0.0004810167, 
    0.0004785863, 0.0004827928, 0.000475234, 0.0004785154, 0.0004725695, 
    0.00047321, 0.0004743689, 0.0004770259, 0.0004755911, 0.0004772689, 
    0.0004735635, 0.000471641, 0.0004711433, 0.0004702151, 0.0004711644, 
    0.0004710871, 0.0004719955, 0.0004717035, 0.0004738844, 0.0004727129, 
    0.0004760406, 0.0004772549, 0.0004806833, 0.0004827847, 0.0004849232, 
    0.0004858673, 0.0004861546, 0.0004862747 ;

 SMINN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_PLANT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_SOIL1N_L1 =
  3.117403e-14, 3.125812e-14, 3.124178e-14, 3.130955e-14, 3.127198e-14, 
    3.131633e-14, 3.11911e-14, 3.126144e-14, 3.121655e-14, 3.118162e-14, 
    3.144085e-14, 3.131257e-14, 3.157399e-14, 3.149233e-14, 3.169734e-14, 
    3.156127e-14, 3.172475e-14, 3.169344e-14, 3.178771e-14, 3.176072e-14, 
    3.18811e-14, 3.180016e-14, 3.194348e-14, 3.186179e-14, 3.187457e-14, 
    3.179749e-14, 3.133843e-14, 3.142488e-14, 3.13333e-14, 3.134563e-14, 
    3.134011e-14, 3.127274e-14, 3.123875e-14, 3.116761e-14, 3.118054e-14, 
    3.12328e-14, 3.135118e-14, 3.131103e-14, 3.141223e-14, 3.140995e-14, 
    3.152244e-14, 3.147174e-14, 3.166058e-14, 3.160698e-14, 3.176184e-14, 
    3.172292e-14, 3.176001e-14, 3.174877e-14, 3.176016e-14, 3.170306e-14, 
    3.172753e-14, 3.167727e-14, 3.148123e-14, 3.15389e-14, 3.136678e-14, 
    3.126307e-14, 3.119418e-14, 3.114524e-14, 3.115216e-14, 3.116534e-14, 
    3.12331e-14, 3.129679e-14, 3.134527e-14, 3.137769e-14, 3.140962e-14, 
    3.150612e-14, 3.155721e-14, 3.167141e-14, 3.165083e-14, 3.168571e-14, 
    3.171904e-14, 3.177495e-14, 3.176575e-14, 3.179037e-14, 3.168481e-14, 
    3.175497e-14, 3.163912e-14, 3.167081e-14, 3.141821e-14, 3.132187e-14, 
    3.128081e-14, 3.124492e-14, 3.115748e-14, 3.121787e-14, 3.119407e-14, 
    3.12507e-14, 3.128666e-14, 3.126889e-14, 3.137858e-14, 3.133595e-14, 
    3.156023e-14, 3.14637e-14, 3.171516e-14, 3.165506e-14, 3.172956e-14, 
    3.169155e-14, 3.175665e-14, 3.169807e-14, 3.179953e-14, 3.18216e-14, 
    3.180652e-14, 3.186446e-14, 3.169482e-14, 3.176e-14, 3.126838e-14, 
    3.127128e-14, 3.12848e-14, 3.122536e-14, 3.122173e-14, 3.116726e-14, 
    3.121574e-14, 3.123637e-14, 3.128875e-14, 3.13197e-14, 3.134912e-14, 
    3.141377e-14, 3.148588e-14, 3.158665e-14, 3.165895e-14, 3.170739e-14, 
    3.16777e-14, 3.170391e-14, 3.167461e-14, 3.166087e-14, 3.181333e-14, 
    3.172775e-14, 3.185613e-14, 3.184904e-14, 3.179095e-14, 3.184984e-14, 
    3.127332e-14, 3.125663e-14, 3.119864e-14, 3.124403e-14, 3.116132e-14, 
    3.120761e-14, 3.123421e-14, 3.133682e-14, 3.135937e-14, 3.138024e-14, 
    3.142147e-14, 3.147434e-14, 3.156699e-14, 3.164752e-14, 3.172099e-14, 
    3.171561e-14, 3.17175e-14, 3.17339e-14, 3.169327e-14, 3.174056e-14, 
    3.174849e-14, 3.172775e-14, 3.184809e-14, 3.181373e-14, 3.184889e-14, 
    3.182652e-14, 3.126206e-14, 3.129014e-14, 3.127496e-14, 3.130349e-14, 
    3.128339e-14, 3.137271e-14, 3.139947e-14, 3.152459e-14, 3.147329e-14, 
    3.155495e-14, 3.14816e-14, 3.14946e-14, 3.155757e-14, 3.148557e-14, 
    3.164306e-14, 3.153629e-14, 3.173453e-14, 3.1628e-14, 3.17412e-14, 
    3.172067e-14, 3.175467e-14, 3.17851e-14, 3.182338e-14, 3.189394e-14, 
    3.187761e-14, 3.19366e-14, 3.133199e-14, 3.136837e-14, 3.136518e-14, 
    3.140325e-14, 3.143139e-14, 3.149236e-14, 3.159003e-14, 3.155332e-14, 
    3.162072e-14, 3.163424e-14, 3.153185e-14, 3.159471e-14, 3.139272e-14, 
    3.142537e-14, 3.140595e-14, 3.133485e-14, 3.156176e-14, 3.144538e-14, 
    3.166015e-14, 3.159722e-14, 3.178076e-14, 3.168951e-14, 3.186862e-14, 
    3.194501e-14, 3.201693e-14, 3.210078e-14, 3.138824e-14, 3.136352e-14, 
    3.140778e-14, 3.146894e-14, 3.15257e-14, 3.160106e-14, 3.160878e-14, 
    3.162288e-14, 3.16594e-14, 3.169011e-14, 3.162732e-14, 3.16978e-14, 
    3.14329e-14, 3.157186e-14, 3.135416e-14, 3.141976e-14, 3.146535e-14, 
    3.144537e-14, 3.154913e-14, 3.157356e-14, 3.167273e-14, 3.16215e-14, 
    3.192615e-14, 3.17915e-14, 3.216462e-14, 3.206053e-14, 3.135488e-14, 
    3.138816e-14, 3.150384e-14, 3.144882e-14, 3.16061e-14, 3.164474e-14, 
    3.167616e-14, 3.171629e-14, 3.172063e-14, 3.17444e-14, 3.170545e-14, 
    3.174287e-14, 3.160122e-14, 3.166454e-14, 3.149064e-14, 3.1533e-14, 
    3.151352e-14, 3.149214e-14, 3.155811e-14, 3.162831e-14, 3.162983e-14, 
    3.16523e-14, 3.171559e-14, 3.160673e-14, 3.194346e-14, 3.173562e-14, 
    3.142442e-14, 3.148841e-14, 3.149758e-14, 3.14728e-14, 3.164088e-14, 
    3.158001e-14, 3.174382e-14, 3.169959e-14, 3.177206e-14, 3.173605e-14, 
    3.173075e-14, 3.168448e-14, 3.165566e-14, 3.15828e-14, 3.152347e-14, 
    3.147639e-14, 3.148735e-14, 3.153904e-14, 3.16326e-14, 3.172101e-14, 
    3.170165e-14, 3.176656e-14, 3.15947e-14, 3.166678e-14, 3.163893e-14, 
    3.171157e-14, 3.155234e-14, 3.168786e-14, 3.151765e-14, 3.153259e-14, 
    3.15788e-14, 3.167165e-14, 3.169223e-14, 3.171414e-14, 3.170062e-14, 
    3.163498e-14, 3.162423e-14, 3.157769e-14, 3.156482e-14, 3.152934e-14, 
    3.149994e-14, 3.15268e-14, 3.155498e-14, 3.163502e-14, 3.170705e-14, 
    3.178553e-14, 3.180474e-14, 3.189624e-14, 3.182172e-14, 3.194461e-14, 
    3.184008e-14, 3.202096e-14, 3.169575e-14, 3.183706e-14, 3.158092e-14, 
    3.160856e-14, 3.165849e-14, 3.177299e-14, 3.171123e-14, 3.178346e-14, 
    3.162381e-14, 3.154081e-14, 3.151936e-14, 3.147925e-14, 3.152027e-14, 
    3.151694e-14, 3.155617e-14, 3.154356e-14, 3.163768e-14, 3.158714e-14, 
    3.173061e-14, 3.17829e-14, 3.193041e-14, 3.202068e-14, 3.21125e-14, 
    3.215298e-14, 3.216531e-14, 3.217045e-14 ;

 SMINN_TO_SOIL1N_L2 =
  1.036534e-14, 1.039333e-14, 1.038789e-14, 1.041044e-14, 1.039794e-14, 
    1.04127e-14, 1.037102e-14, 1.039443e-14, 1.037949e-14, 1.036786e-14, 
    1.045414e-14, 1.041145e-14, 1.049846e-14, 1.047128e-14, 1.053951e-14, 
    1.049422e-14, 1.054863e-14, 1.053821e-14, 1.056959e-14, 1.05606e-14, 
    1.060067e-14, 1.057373e-14, 1.062143e-14, 1.059425e-14, 1.05985e-14, 
    1.057284e-14, 1.042006e-14, 1.044883e-14, 1.041835e-14, 1.042245e-14, 
    1.042061e-14, 1.039819e-14, 1.038688e-14, 1.03632e-14, 1.036751e-14, 
    1.03849e-14, 1.04243e-14, 1.041094e-14, 1.044462e-14, 1.044386e-14, 
    1.04813e-14, 1.046442e-14, 1.052728e-14, 1.050944e-14, 1.056098e-14, 
    1.054802e-14, 1.056037e-14, 1.055663e-14, 1.056042e-14, 1.054141e-14, 
    1.054956e-14, 1.053283e-14, 1.046758e-14, 1.048678e-14, 1.042949e-14, 
    1.039497e-14, 1.037204e-14, 1.035576e-14, 1.035806e-14, 1.036245e-14, 
    1.0385e-14, 1.04062e-14, 1.042233e-14, 1.043312e-14, 1.044375e-14, 
    1.047587e-14, 1.049287e-14, 1.053088e-14, 1.052403e-14, 1.053564e-14, 
    1.054673e-14, 1.056534e-14, 1.056228e-14, 1.057047e-14, 1.053534e-14, 
    1.055869e-14, 1.052013e-14, 1.053068e-14, 1.044661e-14, 1.041454e-14, 
    1.040088e-14, 1.038893e-14, 1.035983e-14, 1.037993e-14, 1.037201e-14, 
    1.039086e-14, 1.040283e-14, 1.039691e-14, 1.043342e-14, 1.041923e-14, 
    1.049388e-14, 1.046175e-14, 1.054544e-14, 1.052544e-14, 1.055023e-14, 
    1.053759e-14, 1.055925e-14, 1.053975e-14, 1.057352e-14, 1.058087e-14, 
    1.057585e-14, 1.059514e-14, 1.053867e-14, 1.056037e-14, 1.039674e-14, 
    1.039771e-14, 1.04022e-14, 1.038243e-14, 1.038122e-14, 1.036308e-14, 
    1.037922e-14, 1.038609e-14, 1.040352e-14, 1.041382e-14, 1.042361e-14, 
    1.044513e-14, 1.046913e-14, 1.050267e-14, 1.052673e-14, 1.054286e-14, 
    1.053297e-14, 1.05417e-14, 1.053194e-14, 1.052737e-14, 1.057812e-14, 
    1.054963e-14, 1.059236e-14, 1.059e-14, 1.057067e-14, 1.059027e-14, 
    1.039838e-14, 1.039283e-14, 1.037353e-14, 1.038864e-14, 1.036111e-14, 
    1.037652e-14, 1.038537e-14, 1.041952e-14, 1.042702e-14, 1.043397e-14, 
    1.044769e-14, 1.046529e-14, 1.049613e-14, 1.052293e-14, 1.054738e-14, 
    1.054559e-14, 1.054622e-14, 1.055168e-14, 1.053815e-14, 1.05539e-14, 
    1.055654e-14, 1.054963e-14, 1.058968e-14, 1.057825e-14, 1.058995e-14, 
    1.058251e-14, 1.039464e-14, 1.040398e-14, 1.039893e-14, 1.040843e-14, 
    1.040174e-14, 1.043146e-14, 1.044037e-14, 1.048202e-14, 1.046494e-14, 
    1.049212e-14, 1.046771e-14, 1.047203e-14, 1.049299e-14, 1.046903e-14, 
    1.052145e-14, 1.048591e-14, 1.055189e-14, 1.051643e-14, 1.055411e-14, 
    1.054728e-14, 1.055859e-14, 1.056872e-14, 1.058146e-14, 1.060495e-14, 
    1.059951e-14, 1.061915e-14, 1.041791e-14, 1.043002e-14, 1.042896e-14, 
    1.044163e-14, 1.045099e-14, 1.047129e-14, 1.050379e-14, 1.049158e-14, 
    1.051401e-14, 1.051851e-14, 1.048443e-14, 1.050535e-14, 1.043812e-14, 
    1.044899e-14, 1.044253e-14, 1.041886e-14, 1.049438e-14, 1.045565e-14, 
    1.052713e-14, 1.050619e-14, 1.056728e-14, 1.05369e-14, 1.059652e-14, 
    1.062194e-14, 1.064588e-14, 1.067379e-14, 1.043663e-14, 1.042841e-14, 
    1.044314e-14, 1.046349e-14, 1.048238e-14, 1.050746e-14, 1.051003e-14, 
    1.051473e-14, 1.052688e-14, 1.05371e-14, 1.051621e-14, 1.053966e-14, 
    1.04515e-14, 1.049775e-14, 1.042529e-14, 1.044712e-14, 1.04623e-14, 
    1.045565e-14, 1.049018e-14, 1.049831e-14, 1.053132e-14, 1.051427e-14, 
    1.061567e-14, 1.057085e-14, 1.069504e-14, 1.066039e-14, 1.042553e-14, 
    1.043661e-14, 1.047511e-14, 1.04568e-14, 1.050914e-14, 1.0522e-14, 
    1.053246e-14, 1.054582e-14, 1.054726e-14, 1.055517e-14, 1.054221e-14, 
    1.055466e-14, 1.050752e-14, 1.052859e-14, 1.047072e-14, 1.048481e-14, 
    1.047833e-14, 1.047121e-14, 1.049317e-14, 1.051653e-14, 1.051704e-14, 
    1.052452e-14, 1.054558e-14, 1.050935e-14, 1.062143e-14, 1.055225e-14, 
    1.044868e-14, 1.046997e-14, 1.047303e-14, 1.046478e-14, 1.052072e-14, 
    1.050046e-14, 1.055498e-14, 1.054026e-14, 1.056438e-14, 1.05524e-14, 
    1.055063e-14, 1.053523e-14, 1.052564e-14, 1.050139e-14, 1.048164e-14, 
    1.046597e-14, 1.046962e-14, 1.048682e-14, 1.051796e-14, 1.054739e-14, 
    1.054094e-14, 1.056255e-14, 1.050535e-14, 1.052934e-14, 1.052007e-14, 
    1.054425e-14, 1.049125e-14, 1.053636e-14, 1.04797e-14, 1.048468e-14, 
    1.050006e-14, 1.053096e-14, 1.053781e-14, 1.05451e-14, 1.05406e-14, 
    1.051876e-14, 1.051518e-14, 1.049969e-14, 1.04954e-14, 1.04836e-14, 
    1.047381e-14, 1.048275e-14, 1.049213e-14, 1.051877e-14, 1.054274e-14, 
    1.056886e-14, 1.057526e-14, 1.060571e-14, 1.058091e-14, 1.062181e-14, 
    1.058702e-14, 1.064722e-14, 1.053898e-14, 1.058602e-14, 1.050076e-14, 
    1.050996e-14, 1.052658e-14, 1.056469e-14, 1.054413e-14, 1.056818e-14, 
    1.051504e-14, 1.048741e-14, 1.048027e-14, 1.046693e-14, 1.048058e-14, 
    1.047947e-14, 1.049252e-14, 1.048833e-14, 1.051965e-14, 1.050283e-14, 
    1.055058e-14, 1.056799e-14, 1.061708e-14, 1.064713e-14, 1.067769e-14, 
    1.069117e-14, 1.069527e-14, 1.069698e-14 ;

 SMINN_TO_SOIL1N_S2 =
  -8.365502e-11, -8.402314e-11, -8.395157e-11, -8.424849e-11, -8.408378e-11, 
    -8.427821e-11, -8.372966e-11, -8.403776e-11, -8.384107e-11, 
    -8.368816e-11, -8.482471e-11, -8.426174e-11, -8.540944e-11, 
    -8.505041e-11, -8.595229e-11, -8.535358e-11, -8.607302e-11, 
    -8.593502e-11, -8.635035e-11, -8.623136e-11, -8.676262e-11, 
    -8.640526e-11, -8.7038e-11, -8.667728e-11, -8.673371e-11, -8.639348e-11, 
    -8.437502e-11, -8.475463e-11, -8.435253e-11, -8.440666e-11, 
    -8.438238e-11, -8.408719e-11, -8.393844e-11, -8.362688e-11, 
    -8.368344e-11, -8.391227e-11, -8.4431e-11, -8.425491e-11, -8.469869e-11, 
    -8.468867e-11, -8.518272e-11, -8.495996e-11, -8.579035e-11, 
    -8.555433e-11, -8.623633e-11, -8.606481e-11, -8.622827e-11, 
    -8.617871e-11, -8.622892e-11, -8.597738e-11, -8.608515e-11, -8.58638e-11, 
    -8.500169e-11, -8.525506e-11, -8.449937e-11, -8.404499e-11, 
    -8.374317e-11, -8.352899e-11, -8.355927e-11, -8.3617e-11, -8.391361e-11, 
    -8.419248e-11, -8.4405e-11, -8.454715e-11, -8.468723e-11, -8.511123e-11, 
    -8.533562e-11, -8.583807e-11, -8.574739e-11, -8.590101e-11, 
    -8.604775e-11, -8.629414e-11, -8.625358e-11, -8.636213e-11, 
    -8.589695e-11, -8.620612e-11, -8.569574e-11, -8.583533e-11, 
    -8.472534e-11, -8.430242e-11, -8.412268e-11, -8.396533e-11, 
    -8.358255e-11, -8.384689e-11, -8.374269e-11, -8.399059e-11, 
    -8.414812e-11, -8.407021e-11, -8.455105e-11, -8.436411e-11, 
    -8.534892e-11, -8.492473e-11, -8.603063e-11, -8.5766e-11, -8.609406e-11, 
    -8.592666e-11, -8.62135e-11, -8.595535e-11, -8.640253e-11, -8.649991e-11, 
    -8.643337e-11, -8.668898e-11, -8.594104e-11, -8.622827e-11, 
    -8.406803e-11, -8.408074e-11, -8.413993e-11, -8.387972e-11, -8.38638e-11, 
    -8.362533e-11, -8.383752e-11, -8.392788e-11, -8.415725e-11, 
    -8.429293e-11, -8.44219e-11, -8.470547e-11, -8.502217e-11, -8.546502e-11, 
    -8.578315e-11, -8.599641e-11, -8.586564e-11, -8.59811e-11, -8.585203e-11, 
    -8.579154e-11, -8.646343e-11, -8.608616e-11, -8.665221e-11, 
    -8.662088e-11, -8.636472e-11, -8.662442e-11, -8.408966e-11, 
    -8.401654e-11, -8.376267e-11, -8.396134e-11, -8.359936e-11, 
    -8.380199e-11, -8.39185e-11, -8.436803e-11, -8.446678e-11, -8.455837e-11, 
    -8.473924e-11, -8.497136e-11, -8.537857e-11, -8.573287e-11, 
    -8.605629e-11, -8.603259e-11, -8.604093e-11, -8.611319e-11, 
    -8.593422e-11, -8.614257e-11, -8.617754e-11, -8.608611e-11, 
    -8.661669e-11, -8.646511e-11, -8.662022e-11, -8.652152e-11, -8.40403e-11, 
    -8.416334e-11, -8.409685e-11, -8.422188e-11, -8.41338e-11, -8.452545e-11, 
    -8.464287e-11, -8.519229e-11, -8.49668e-11, -8.532566e-11, -8.500325e-11, 
    -8.506038e-11, -8.533739e-11, -8.502067e-11, -8.571334e-11, 
    -8.524374e-11, -8.6116e-11, -8.564708e-11, -8.614538e-11, -8.605489e-11, 
    -8.620471e-11, -8.63389e-11, -8.650771e-11, -8.68192e-11, -8.674707e-11, 
    -8.700755e-11, -8.434676e-11, -8.450635e-11, -8.449229e-11, 
    -8.465929e-11, -8.478281e-11, -8.505049e-11, -8.547984e-11, 
    -8.531838e-11, -8.561479e-11, -8.567429e-11, -8.522399e-11, 
    -8.550047e-11, -8.461315e-11, -8.475651e-11, -8.467115e-11, 
    -8.435935e-11, -8.53556e-11, -8.484433e-11, -8.578841e-11, -8.551145e-11, 
    -8.631977e-11, -8.591778e-11, -8.670736e-11, -8.704491e-11, 
    -8.736258e-11, -8.773383e-11, -8.459344e-11, -8.4485e-11, -8.467915e-11, 
    -8.494778e-11, -8.5197e-11, -8.552834e-11, -8.556224e-11, -8.562431e-11, 
    -8.578509e-11, -8.592028e-11, -8.564395e-11, -8.595417e-11, 
    -8.478978e-11, -8.539998e-11, -8.444401e-11, -8.473189e-11, 
    -8.493194e-11, -8.484417e-11, -8.529993e-11, -8.540735e-11, 
    -8.584386e-11, -8.561821e-11, -8.696161e-11, -8.636725e-11, 
    -8.801649e-11, -8.755561e-11, -8.444712e-11, -8.459306e-11, -8.5101e-11, 
    -8.485932e-11, -8.555046e-11, -8.572058e-11, -8.585887e-11, 
    -8.603566e-11, -8.605474e-11, -8.615949e-11, -8.598784e-11, 
    -8.615271e-11, -8.552905e-11, -8.580774e-11, -8.504293e-11, 
    -8.522909e-11, -8.514345e-11, -8.504951e-11, -8.533942e-11, -8.56483e-11, 
    -8.565489e-11, -8.575393e-11, -8.603305e-11, -8.555326e-11, 
    -8.703834e-11, -8.612121e-11, -8.475221e-11, -8.503333e-11, 
    -8.507347e-11, -8.496457e-11, -8.570353e-11, -8.543578e-11, 
    -8.615694e-11, -8.596203e-11, -8.628138e-11, -8.612269e-11, 
    -8.609934e-11, -8.589553e-11, -8.576864e-11, -8.544806e-11, 
    -8.518721e-11, -8.498036e-11, -8.502846e-11, -8.525568e-11, 
    -8.566719e-11, -8.605647e-11, -8.59712e-11, -8.625711e-11, -8.550034e-11, 
    -8.581767e-11, -8.569503e-11, -8.601482e-11, -8.53141e-11, -8.591083e-11, 
    -8.516157e-11, -8.522726e-11, -8.543046e-11, -8.58392e-11, -8.592962e-11, 
    -8.602618e-11, -8.596659e-11, -8.567764e-11, -8.563029e-11, 
    -8.542552e-11, -8.536899e-11, -8.521296e-11, -8.508379e-11, 
    -8.520181e-11, -8.532576e-11, -8.567776e-11, -8.599497e-11, 
    -8.634081e-11, -8.642544e-11, -8.682956e-11, -8.650061e-11, 
    -8.704346e-11, -8.658196e-11, -8.738082e-11, -8.59454e-11, -8.656836e-11, 
    -8.54397e-11, -8.556129e-11, -8.578123e-11, -8.628565e-11, -8.601331e-11, 
    -8.63318e-11, -8.562843e-11, -8.526353e-11, -8.516909e-11, -8.499294e-11, 
    -8.517313e-11, -8.515846e-11, -8.533088e-11, -8.527547e-11, 
    -8.568944e-11, -8.546708e-11, -8.609876e-11, -8.632928e-11, 
    -8.698026e-11, -8.737933e-11, -8.778554e-11, -8.796489e-11, 
    -8.801947e-11, -8.804229e-11 ;

 SMINN_TO_SOIL1N_S3 =
  -2.016235e-12, -2.025105e-12, -2.023381e-12, -2.030535e-12, -2.026566e-12, 
    -2.031251e-12, -2.018033e-12, -2.025457e-12, -2.020718e-12, 
    -2.017033e-12, -2.04442e-12, -2.030854e-12, -2.05851e-12, -2.049858e-12, 
    -2.071591e-12, -2.057164e-12, -2.074499e-12, -2.071174e-12, 
    -2.081182e-12, -2.078315e-12, -2.091116e-12, -2.082505e-12, 
    -2.097752e-12, -2.08906e-12, -2.09042e-12, -2.082221e-12, -2.033584e-12, 
    -2.042731e-12, -2.033042e-12, -2.034346e-12, -2.033761e-12, 
    -2.026648e-12, -2.023064e-12, -2.015557e-12, -2.016919e-12, 
    -2.022433e-12, -2.034933e-12, -2.03069e-12, -2.041383e-12, -2.041142e-12, 
    -2.053047e-12, -2.047679e-12, -2.067688e-12, -2.062001e-12, 
    -2.078435e-12, -2.074302e-12, -2.078241e-12, -2.077046e-12, 
    -2.078256e-12, -2.072195e-12, -2.074792e-12, -2.069458e-12, 
    -2.048684e-12, -2.05479e-12, -2.036581e-12, -2.025632e-12, -2.018359e-12, 
    -2.013198e-12, -2.013927e-12, -2.015318e-12, -2.022466e-12, 
    -2.029185e-12, -2.034306e-12, -2.037732e-12, -2.041107e-12, 
    -2.051324e-12, -2.056731e-12, -2.068838e-12, -2.066653e-12, 
    -2.070355e-12, -2.073891e-12, -2.079828e-12, -2.07885e-12, -2.081466e-12, 
    -2.070257e-12, -2.077707e-12, -2.065408e-12, -2.068772e-12, 
    -2.042026e-12, -2.031835e-12, -2.027504e-12, -2.023712e-12, 
    -2.014488e-12, -2.020858e-12, -2.018347e-12, -2.024321e-12, 
    -2.028117e-12, -2.026239e-12, -2.037826e-12, -2.033321e-12, 
    -2.057052e-12, -2.04683e-12, -2.073478e-12, -2.067101e-12, -2.075007e-12, 
    -2.070973e-12, -2.077885e-12, -2.071664e-12, -2.082439e-12, 
    -2.084786e-12, -2.083183e-12, -2.089342e-12, -2.071319e-12, 
    -2.078241e-12, -2.026187e-12, -2.026493e-12, -2.027919e-12, 
    -2.021649e-12, -2.021266e-12, -2.015519e-12, -2.020632e-12, 
    -2.022809e-12, -2.028336e-12, -2.031606e-12, -2.034714e-12, 
    -2.041547e-12, -2.049178e-12, -2.059849e-12, -2.067515e-12, 
    -2.072654e-12, -2.069503e-12, -2.072284e-12, -2.069175e-12, 
    -2.067717e-12, -2.083907e-12, -2.074816e-12, -2.088456e-12, 
    -2.087701e-12, -2.081528e-12, -2.087786e-12, -2.026708e-12, 
    -2.024946e-12, -2.018828e-12, -2.023616e-12, -2.014893e-12, 
    -2.019776e-12, -2.022583e-12, -2.033416e-12, -2.035795e-12, 
    -2.038002e-12, -2.04236e-12, -2.047954e-12, -2.057766e-12, -2.066303e-12, 
    -2.074096e-12, -2.073525e-12, -2.073726e-12, -2.075467e-12, 
    -2.071155e-12, -2.076175e-12, -2.077018e-12, -2.074815e-12, -2.0876e-12, 
    -2.083947e-12, -2.087685e-12, -2.085307e-12, -2.025518e-12, 
    -2.028483e-12, -2.026881e-12, -2.029894e-12, -2.027771e-12, 
    -2.037209e-12, -2.040038e-12, -2.053277e-12, -2.047844e-12, 
    -2.056491e-12, -2.048722e-12, -2.050099e-12, -2.056774e-12, 
    -2.049142e-12, -2.065833e-12, -2.054517e-12, -2.075535e-12, 
    -2.064236e-12, -2.076243e-12, -2.074063e-12, -2.077673e-12, 
    -2.080906e-12, -2.084974e-12, -2.09248e-12, -2.090741e-12, -2.097018e-12, 
    -2.032903e-12, -2.036749e-12, -2.03641e-12, -2.040434e-12, -2.04341e-12, 
    -2.04986e-12, -2.060206e-12, -2.056316e-12, -2.063458e-12, -2.064892e-12, 
    -2.054041e-12, -2.060703e-12, -2.039322e-12, -2.042777e-12, -2.04072e-12, 
    -2.033207e-12, -2.057212e-12, -2.044893e-12, -2.067642e-12, 
    -2.060968e-12, -2.080445e-12, -2.070759e-12, -2.089785e-12, 
    -2.097918e-12, -2.105573e-12, -2.114519e-12, -2.038847e-12, 
    -2.036234e-12, -2.040913e-12, -2.047385e-12, -2.053391e-12, 
    -2.061375e-12, -2.062192e-12, -2.063687e-12, -2.067562e-12, 
    -2.070819e-12, -2.06416e-12, -2.071636e-12, -2.043578e-12, -2.058282e-12, 
    -2.035246e-12, -2.042183e-12, -2.047004e-12, -2.044889e-12, 
    -2.055871e-12, -2.058459e-12, -2.068978e-12, -2.06354e-12, -2.095911e-12, 
    -2.081589e-12, -2.12133e-12, -2.110224e-12, -2.035321e-12, -2.038838e-12, 
    -2.051077e-12, -2.045254e-12, -2.061908e-12, -2.066007e-12, 
    -2.069339e-12, -2.073599e-12, -2.074059e-12, -2.076583e-12, 
    -2.072447e-12, -2.07642e-12, -2.061392e-12, -2.068107e-12, -2.049678e-12, 
    -2.054164e-12, -2.0521e-12, -2.049837e-12, -2.056823e-12, -2.064265e-12, 
    -2.064424e-12, -2.066811e-12, -2.073536e-12, -2.061975e-12, -2.09776e-12, 
    -2.075661e-12, -2.042673e-12, -2.049447e-12, -2.050414e-12, -2.04779e-12, 
    -2.065596e-12, -2.059144e-12, -2.076521e-12, -2.071825e-12, -2.07952e-12, 
    -2.075696e-12, -2.075134e-12, -2.070223e-12, -2.067165e-12, -2.05944e-12, 
    -2.053155e-12, -2.04817e-12, -2.049329e-12, -2.054805e-12, -2.064721e-12, 
    -2.074101e-12, -2.072046e-12, -2.078935e-12, -2.0607e-12, -2.068347e-12, 
    -2.065391e-12, -2.073097e-12, -2.056212e-12, -2.070592e-12, 
    -2.052537e-12, -2.05412e-12, -2.059016e-12, -2.068865e-12, -2.071044e-12, 
    -2.073371e-12, -2.071935e-12, -2.064972e-12, -2.063831e-12, 
    -2.058897e-12, -2.057535e-12, -2.053775e-12, -2.050663e-12, 
    -2.053507e-12, -2.056493e-12, -2.064975e-12, -2.072619e-12, 
    -2.080952e-12, -2.082992e-12, -2.092729e-12, -2.084803e-12, 
    -2.097883e-12, -2.086763e-12, -2.106012e-12, -2.071424e-12, 
    -2.086435e-12, -2.059239e-12, -2.062169e-12, -2.067468e-12, 
    -2.079623e-12, -2.073061e-12, -2.080735e-12, -2.063787e-12, 
    -2.054994e-12, -2.052718e-12, -2.048474e-12, -2.052815e-12, 
    -2.052462e-12, -2.056617e-12, -2.055282e-12, -2.065257e-12, 
    -2.059898e-12, -2.07512e-12, -2.080674e-12, -2.09636e-12, -2.105977e-12, 
    -2.115765e-12, -2.120086e-12, -2.121401e-12, -2.121951e-12 ;

 SMINN_TO_SOIL2N_L3 =
  3.367222e-15, 3.376314e-15, 3.374547e-15, 3.381874e-15, 3.377812e-15, 
    3.382607e-15, 3.369067e-15, 3.376673e-15, 3.371819e-15, 3.368042e-15, 
    3.39607e-15, 3.382201e-15, 3.410466e-15, 3.401636e-15, 3.423802e-15, 
    3.40909e-15, 3.426766e-15, 3.423381e-15, 3.433573e-15, 3.430655e-15, 
    3.443671e-15, 3.43492e-15, 3.450415e-15, 3.441583e-15, 3.442964e-15, 
    3.43463e-15, 3.384996e-15, 3.394344e-15, 3.384442e-15, 3.385776e-15, 
    3.385178e-15, 3.377895e-15, 3.37422e-15, 3.366528e-15, 3.367926e-15, 
    3.373576e-15, 3.386375e-15, 3.382034e-15, 3.392976e-15, 3.392729e-15, 
    3.404892e-15, 3.39941e-15, 3.419828e-15, 3.414032e-15, 3.430776e-15, 
    3.426567e-15, 3.430578e-15, 3.429363e-15, 3.430594e-15, 3.424421e-15, 
    3.427066e-15, 3.421633e-15, 3.400437e-15, 3.406671e-15, 3.388062e-15, 
    3.376849e-15, 3.3694e-15, 3.364109e-15, 3.364857e-15, 3.366283e-15, 
    3.373609e-15, 3.380494e-15, 3.385737e-15, 3.389241e-15, 3.392694e-15, 
    3.403127e-15, 3.40865e-15, 3.420999e-15, 3.418774e-15, 3.422544e-15, 
    3.426149e-15, 3.432193e-15, 3.431199e-15, 3.433861e-15, 3.422447e-15, 
    3.430033e-15, 3.417507e-15, 3.420933e-15, 3.393622e-15, 3.383206e-15, 
    3.378767e-15, 3.374887e-15, 3.365432e-15, 3.371962e-15, 3.369388e-15, 
    3.375512e-15, 3.3794e-15, 3.377477e-15, 3.389337e-15, 3.384728e-15, 
    3.408978e-15, 3.398541e-15, 3.425728e-15, 3.419231e-15, 3.427286e-15, 
    3.423177e-15, 3.430215e-15, 3.423881e-15, 3.434852e-15, 3.437237e-15, 
    3.435607e-15, 3.441872e-15, 3.423529e-15, 3.430577e-15, 3.377423e-15, 
    3.377737e-15, 3.379198e-15, 3.372772e-15, 3.37238e-15, 3.366489e-15, 
    3.371732e-15, 3.373962e-15, 3.379626e-15, 3.382972e-15, 3.386153e-15, 
    3.393142e-15, 3.400939e-15, 3.411834e-15, 3.419652e-15, 3.424889e-15, 
    3.421679e-15, 3.424513e-15, 3.421344e-15, 3.419859e-15, 3.436343e-15, 
    3.42709e-15, 3.440971e-15, 3.440204e-15, 3.433923e-15, 3.440291e-15, 
    3.377957e-15, 3.376153e-15, 3.369882e-15, 3.37479e-15, 3.365848e-15, 
    3.370853e-15, 3.373729e-15, 3.384822e-15, 3.38726e-15, 3.389517e-15, 
    3.393975e-15, 3.399691e-15, 3.409709e-15, 3.418415e-15, 3.426359e-15, 
    3.425777e-15, 3.425982e-15, 3.427755e-15, 3.423362e-15, 3.428476e-15, 
    3.429333e-15, 3.42709e-15, 3.440101e-15, 3.436386e-15, 3.440188e-15, 
    3.437769e-15, 3.376739e-15, 3.379775e-15, 3.378135e-15, 3.381219e-15, 
    3.379045e-15, 3.388703e-15, 3.391596e-15, 3.405125e-15, 3.399578e-15, 
    3.408407e-15, 3.400476e-15, 3.401881e-15, 3.408691e-15, 3.400905e-15, 
    3.417933e-15, 3.406389e-15, 3.427823e-15, 3.416305e-15, 3.428545e-15, 
    3.426325e-15, 3.430001e-15, 3.433291e-15, 3.43743e-15, 3.445059e-15, 
    3.443294e-15, 3.449672e-15, 3.3843e-15, 3.388233e-15, 3.387889e-15, 
    3.392005e-15, 3.395047e-15, 3.401639e-15, 3.4122e-15, 3.408231e-15, 
    3.415518e-15, 3.416979e-15, 3.405909e-15, 3.412706e-15, 3.390866e-15, 
    3.394396e-15, 3.392296e-15, 3.384609e-15, 3.409143e-15, 3.39656e-15, 
    3.419781e-15, 3.412977e-15, 3.432822e-15, 3.422955e-15, 3.442321e-15, 
    3.450581e-15, 3.458357e-15, 3.467423e-15, 3.390381e-15, 3.387709e-15, 
    3.392495e-15, 3.399107e-15, 3.405244e-15, 3.413392e-15, 3.414226e-15, 
    3.415751e-15, 3.4197e-15, 3.42302e-15, 3.416231e-15, 3.423852e-15, 
    3.395211e-15, 3.410235e-15, 3.386697e-15, 3.393789e-15, 3.398719e-15, 
    3.396558e-15, 3.407777e-15, 3.410419e-15, 3.421141e-15, 3.415602e-15, 
    3.448542e-15, 3.433983e-15, 3.474326e-15, 3.46307e-15, 3.386775e-15, 
    3.390373e-15, 3.40288e-15, 3.396932e-15, 3.413937e-15, 3.418114e-15, 
    3.421512e-15, 3.425851e-15, 3.42632e-15, 3.42889e-15, 3.424679e-15, 
    3.428725e-15, 3.413409e-15, 3.420256e-15, 3.401454e-15, 3.406033e-15, 
    3.403927e-15, 3.401615e-15, 3.408748e-15, 3.416338e-15, 3.416503e-15, 
    3.418933e-15, 3.425775e-15, 3.414005e-15, 3.450413e-15, 3.427941e-15, 
    3.394294e-15, 3.401213e-15, 3.402204e-15, 3.399524e-15, 3.417697e-15, 
    3.411117e-15, 3.428828e-15, 3.424045e-15, 3.431881e-15, 3.427988e-15, 
    3.427415e-15, 3.422412e-15, 3.419295e-15, 3.411418e-15, 3.405003e-15, 
    3.399913e-15, 3.401097e-15, 3.406687e-15, 3.416803e-15, 3.426362e-15, 
    3.424268e-15, 3.431286e-15, 3.412705e-15, 3.420498e-15, 3.417487e-15, 
    3.42534e-15, 3.408124e-15, 3.422777e-15, 3.404373e-15, 3.405989e-15, 
    3.410986e-15, 3.421025e-15, 3.423249e-15, 3.425618e-15, 3.424157e-15, 
    3.41706e-15, 3.415898e-15, 3.410865e-15, 3.409474e-15, 3.405638e-15, 
    3.402459e-15, 3.405363e-15, 3.40841e-15, 3.417064e-15, 3.424852e-15, 
    3.433338e-15, 3.435414e-15, 3.445307e-15, 3.43725e-15, 3.450537e-15, 
    3.439235e-15, 3.458793e-15, 3.42363e-15, 3.43891e-15, 3.411214e-15, 
    3.414203e-15, 3.419602e-15, 3.431981e-15, 3.425303e-15, 3.433114e-15, 
    3.415852e-15, 3.406878e-15, 3.404558e-15, 3.400222e-15, 3.404657e-15, 
    3.404297e-15, 3.408539e-15, 3.407176e-15, 3.417351e-15, 3.411887e-15, 
    3.4274e-15, 3.433053e-15, 3.449002e-15, 3.458762e-15, 3.46869e-15, 
    3.473068e-15, 3.4744e-15, 3.474956e-15 ;

 SMINN_TO_SOIL2N_S1 =
  -8.758231e-09, -8.796739e-09, -8.789253e-09, -8.820313e-09, -8.803083e-09, 
    -8.823421e-09, -8.766038e-09, -8.798269e-09, -8.777693e-09, 
    -8.761697e-09, -8.88059e-09, -8.821699e-09, -8.941757e-09, -8.9042e-09, 
    -8.998543e-09, -8.935913e-09, -9.011171e-09, -8.996735e-09, 
    -9.040182e-09, -9.027735e-09, -9.083308e-09, -9.045927e-09, 
    -9.112114e-09, -9.07438e-09, -9.080283e-09, -9.044694e-09, -8.833549e-09, 
    -8.873259e-09, -8.831196e-09, -8.836859e-09, -8.834318e-09, 
    -8.803439e-09, -8.787879e-09, -8.755287e-09, -8.761203e-09, 
    -8.785142e-09, -8.839406e-09, -8.820985e-09, -8.867407e-09, 
    -8.866359e-09, -8.918041e-09, -8.894738e-09, -8.981602e-09, 
    -8.956914e-09, -9.028255e-09, -9.010313e-09, -9.027412e-09, 
    -9.022227e-09, -9.02748e-09, -9.001167e-09, -9.012441e-09, -8.989287e-09, 
    -8.899103e-09, -8.925608e-09, -8.846557e-09, -8.799026e-09, 
    -8.767452e-09, -8.745046e-09, -8.748215e-09, -8.754252e-09, 
    -8.785281e-09, -8.814453e-09, -8.836684e-09, -8.851556e-09, 
    -8.866208e-09, -8.910562e-09, -8.934036e-09, -8.986595e-09, 
    -8.977109e-09, -8.993178e-09, -9.008528e-09, -9.034302e-09, 
    -9.030059e-09, -9.041415e-09, -8.992753e-09, -9.025094e-09, 
    -8.971706e-09, -8.986308e-09, -8.870195e-09, -8.825954e-09, 
    -8.807152e-09, -8.790693e-09, -8.75065e-09, -8.778303e-09, -8.767402e-09, 
    -8.793335e-09, -8.809813e-09, -8.801663e-09, -8.851963e-09, 
    -8.832408e-09, -8.935427e-09, -8.891053e-09, -9.006738e-09, 
    -8.979056e-09, -9.013373e-09, -8.995862e-09, -9.025867e-09, 
    -8.998862e-09, -9.045641e-09, -9.055827e-09, -9.048866e-09, 
    -9.075604e-09, -8.997366e-09, -9.027413e-09, -8.801435e-09, 
    -8.802764e-09, -8.808956e-09, -8.781736e-09, -8.780071e-09, 
    -8.755125e-09, -8.777322e-09, -8.786774e-09, -8.810768e-09, 
    -8.824961e-09, -8.838453e-09, -8.868117e-09, -8.901246e-09, 
    -8.947571e-09, -8.98085e-09, -9.003158e-09, -8.989478e-09, -9.001556e-09, 
    -8.988056e-09, -8.981727e-09, -9.052011e-09, -9.012546e-09, 
    -9.071758e-09, -9.068482e-09, -9.041685e-09, -9.068851e-09, 
    -8.803697e-09, -8.796048e-09, -8.769492e-09, -8.790274e-09, 
    -8.752408e-09, -8.773604e-09, -8.785793e-09, -8.832817e-09, 
    -8.843148e-09, -8.852728e-09, -8.871649e-09, -8.895931e-09, 
    -8.938528e-09, -8.975589e-09, -9.009422e-09, -9.006943e-09, 
    -9.007815e-09, -9.015373e-09, -8.996651e-09, -9.018447e-09, 
    -9.022106e-09, -9.012541e-09, -9.068043e-09, -9.052187e-09, 
    -9.068412e-09, -9.058088e-09, -8.798534e-09, -8.811405e-09, 
    -8.804451e-09, -8.817529e-09, -8.808315e-09, -8.849285e-09, 
    -8.861567e-09, -8.919042e-09, -8.895453e-09, -8.932994e-09, 
    -8.899266e-09, -8.905243e-09, -8.93422e-09, -8.901089e-09, -8.973546e-09, 
    -8.924424e-09, -9.015667e-09, -8.966616e-09, -9.018741e-09, 
    -9.009275e-09, -9.024948e-09, -9.038985e-09, -9.056643e-09, 
    -9.089226e-09, -9.08168e-09, -9.108929e-09, -8.830592e-09, -8.847286e-09, 
    -8.845817e-09, -8.863286e-09, -8.876206e-09, -8.904209e-09, 
    -8.949121e-09, -8.932232e-09, -8.963237e-09, -8.969462e-09, 
    -8.922357e-09, -8.95128e-09, -8.858459e-09, -8.873457e-09, -8.864526e-09, 
    -8.831909e-09, -8.936125e-09, -8.882642e-09, -8.981401e-09, 
    -8.952427e-09, -9.036983e-09, -8.994933e-09, -9.077527e-09, 
    -9.112838e-09, -9.146065e-09, -9.184901e-09, -8.856397e-09, 
    -8.845054e-09, -8.865364e-09, -8.893464e-09, -8.919534e-09, 
    -8.954195e-09, -8.957741e-09, -8.964235e-09, -8.981053e-09, 
    -8.995194e-09, -8.966288e-09, -8.99874e-09, -8.876936e-09, -8.940767e-09, 
    -8.840765e-09, -8.87088e-09, -8.891807e-09, -8.882626e-09, -8.930302e-09, 
    -8.941538e-09, -8.987199e-09, -8.963595e-09, -9.104123e-09, -9.04195e-09, 
    -9.214468e-09, -9.166258e-09, -8.841091e-09, -8.856357e-09, 
    -8.909492e-09, -8.884211e-09, -8.956508e-09, -8.974304e-09, 
    -8.988771e-09, -9.007263e-09, -9.00926e-09, -9.020217e-09, -9.002262e-09, 
    -9.019508e-09, -8.954268e-09, -8.983422e-09, -8.903418e-09, 
    -8.922891e-09, -8.913932e-09, -8.904106e-09, -8.934433e-09, 
    -8.966744e-09, -8.967433e-09, -8.977793e-09, -9.006991e-09, 
    -8.956802e-09, -9.11215e-09, -9.016213e-09, -8.873005e-09, -8.902413e-09, 
    -8.906611e-09, -8.895221e-09, -8.972521e-09, -8.944512e-09, -9.01995e-09, 
    -8.999561e-09, -9.032967e-09, -9.016367e-09, -9.013925e-09, 
    -8.992605e-09, -8.979331e-09, -8.945796e-09, -8.91851e-09, -8.896873e-09, 
    -8.901903e-09, -8.925673e-09, -8.96872e-09, -9.009441e-09, -9.000521e-09, 
    -9.030428e-09, -8.951266e-09, -8.984461e-09, -8.971631e-09, 
    -9.005084e-09, -8.931783e-09, -8.994206e-09, -8.915828e-09, -8.9227e-09, 
    -8.943956e-09, -8.986714e-09, -8.996171e-09, -9.006272e-09, 
    -9.000039e-09, -8.969812e-09, -8.964859e-09, -8.943439e-09, 
    -8.937525e-09, -8.921203e-09, -8.907691e-09, -8.920037e-09, 
    -8.933003e-09, -8.969824e-09, -9.003007e-09, -9.039185e-09, 
    -9.048037e-09, -9.09031e-09, -9.0559e-09, -9.112684e-09, -9.06441e-09, 
    -9.147975e-09, -8.997822e-09, -9.062988e-09, -8.944923e-09, 
    -8.957642e-09, -8.980648e-09, -9.033413e-09, -9.004927e-09, 
    -9.038241e-09, -8.964665e-09, -8.926493e-09, -8.916615e-09, 
    -8.898188e-09, -8.917037e-09, -8.915503e-09, -8.933539e-09, 
    -8.927744e-09, -8.971047e-09, -8.947787e-09, -9.013864e-09, 
    -9.037977e-09, -9.106073e-09, -9.147819e-09, -9.19031e-09, -9.20907e-09, 
    -9.21478e-09, -9.217167e-09 ;

 SMINN_TO_SOIL3N_S1 =
  -1.039262e-10, -1.043833e-10, -1.042944e-10, -1.046631e-10, -1.044586e-10, 
    -1.047e-10, -1.040189e-10, -1.044015e-10, -1.041572e-10, -1.039673e-10, 
    -1.053787e-10, -1.046796e-10, -1.061048e-10, -1.05659e-10, -1.067789e-10, 
    -1.060354e-10, -1.069288e-10, -1.067575e-10, -1.072732e-10, 
    -1.071255e-10, -1.077852e-10, -1.073414e-10, -1.081272e-10, 
    -1.076792e-10, -1.077493e-10, -1.073268e-10, -1.048203e-10, 
    -1.052917e-10, -1.047923e-10, -1.048596e-10, -1.048294e-10, 
    -1.044628e-10, -1.042781e-10, -1.038912e-10, -1.039615e-10, 
    -1.042456e-10, -1.048898e-10, -1.046711e-10, -1.052222e-10, 
    -1.052098e-10, -1.058233e-10, -1.055466e-10, -1.065778e-10, 
    -1.062847e-10, -1.071316e-10, -1.069187e-10, -1.071216e-10, 
    -1.070601e-10, -1.071224e-10, -1.068101e-10, -1.069439e-10, -1.06669e-10, 
    -1.055985e-10, -1.059131e-10, -1.049747e-10, -1.044104e-10, 
    -1.040356e-10, -1.037697e-10, -1.038073e-10, -1.03879e-10, -1.042473e-10, 
    -1.045936e-10, -1.048575e-10, -1.05034e-10, -1.05208e-10, -1.057345e-10, 
    -1.060131e-10, -1.066371e-10, -1.065245e-10, -1.067152e-10, 
    -1.068975e-10, -1.072034e-10, -1.071531e-10, -1.072879e-10, 
    -1.067102e-10, -1.070941e-10, -1.064603e-10, -1.066337e-10, 
    -1.052553e-10, -1.047301e-10, -1.045069e-10, -1.043115e-10, 
    -1.038362e-10, -1.041645e-10, -1.040351e-10, -1.043429e-10, 
    -1.045385e-10, -1.044418e-10, -1.050389e-10, -1.048067e-10, 
    -1.060297e-10, -1.055029e-10, -1.068762e-10, -1.065476e-10, -1.06955e-10, 
    -1.067471e-10, -1.071033e-10, -1.067827e-10, -1.07338e-10, -1.07459e-10, 
    -1.073763e-10, -1.076937e-10, -1.067649e-10, -1.071216e-10, -1.04439e-10, 
    -1.044548e-10, -1.045283e-10, -1.042052e-10, -1.041854e-10, 
    -1.038893e-10, -1.041528e-10, -1.04265e-10, -1.045498e-10, -1.047183e-10, 
    -1.048785e-10, -1.052306e-10, -1.056239e-10, -1.061738e-10, 
    -1.065689e-10, -1.068337e-10, -1.066713e-10, -1.068147e-10, 
    -1.066544e-10, -1.065793e-10, -1.074137e-10, -1.069452e-10, 
    -1.076481e-10, -1.076092e-10, -1.072911e-10, -1.076136e-10, 
    -1.044659e-10, -1.043751e-10, -1.040599e-10, -1.043066e-10, 
    -1.038571e-10, -1.041087e-10, -1.042534e-10, -1.048116e-10, 
    -1.049342e-10, -1.050479e-10, -1.052725e-10, -1.055608e-10, 
    -1.060665e-10, -1.065064e-10, -1.069081e-10, -1.068786e-10, -1.06889e-10, 
    -1.069787e-10, -1.067565e-10, -1.070152e-10, -1.070586e-10, 
    -1.069451e-10, -1.07604e-10, -1.074157e-10, -1.076084e-10, -1.074858e-10, 
    -1.044046e-10, -1.045574e-10, -1.044748e-10, -1.046301e-10, 
    -1.045207e-10, -1.050071e-10, -1.051529e-10, -1.058351e-10, 
    -1.055551e-10, -1.060008e-10, -1.056004e-10, -1.056713e-10, 
    -1.060153e-10, -1.05622e-10, -1.064822e-10, -1.05899e-10, -1.069822e-10, 
    -1.063999e-10, -1.070187e-10, -1.069063e-10, -1.070924e-10, -1.07259e-10, 
    -1.074686e-10, -1.078555e-10, -1.077659e-10, -1.080894e-10, 
    -1.047852e-10, -1.049833e-10, -1.049659e-10, -1.051733e-10, 
    -1.053266e-10, -1.056591e-10, -1.061922e-10, -1.059917e-10, 
    -1.063598e-10, -1.064337e-10, -1.058745e-10, -1.062178e-10, -1.05116e-10, 
    -1.05294e-10, -1.05188e-10, -1.048008e-10, -1.060379e-10, -1.05403e-10, 
    -1.065754e-10, -1.062315e-10, -1.072353e-10, -1.067361e-10, 
    -1.077166e-10, -1.081358e-10, -1.085303e-10, -1.089913e-10, 
    -1.050915e-10, -1.049568e-10, -1.051979e-10, -1.055315e-10, -1.05841e-10, 
    -1.062525e-10, -1.062945e-10, -1.063716e-10, -1.065713e-10, 
    -1.067392e-10, -1.06396e-10, -1.067813e-10, -1.053353e-10, -1.060931e-10, 
    -1.049059e-10, -1.052634e-10, -1.055118e-10, -1.054029e-10, 
    -1.059688e-10, -1.061022e-10, -1.066443e-10, -1.06364e-10, -1.080323e-10, 
    -1.072942e-10, -1.093423e-10, -1.0877e-10, -1.049098e-10, -1.05091e-10, 
    -1.057218e-10, -1.054217e-10, -1.062799e-10, -1.064912e-10, 
    -1.066629e-10, -1.068824e-10, -1.069061e-10, -1.070362e-10, 
    -1.068231e-10, -1.070278e-10, -1.062533e-10, -1.065994e-10, 
    -1.056497e-10, -1.058808e-10, -1.057745e-10, -1.056578e-10, 
    -1.060179e-10, -1.064014e-10, -1.064096e-10, -1.065326e-10, 
    -1.068792e-10, -1.062834e-10, -1.081276e-10, -1.069887e-10, 
    -1.052886e-10, -1.056377e-10, -1.056876e-10, -1.055524e-10, -1.0647e-10, 
    -1.061375e-10, -1.07033e-10, -1.06791e-10, -1.071876e-10, -1.069905e-10, 
    -1.069615e-10, -1.067084e-10, -1.065509e-10, -1.061528e-10, 
    -1.058288e-10, -1.05572e-10, -1.056317e-10, -1.059139e-10, -1.064249e-10, 
    -1.069083e-10, -1.068024e-10, -1.071574e-10, -1.062177e-10, 
    -1.066117e-10, -1.064595e-10, -1.068566e-10, -1.059864e-10, 
    -1.067274e-10, -1.05797e-10, -1.058786e-10, -1.061309e-10, -1.066385e-10, 
    -1.067508e-10, -1.068707e-10, -1.067967e-10, -1.064379e-10, 
    -1.063791e-10, -1.061248e-10, -1.060546e-10, -1.058608e-10, 
    -1.057004e-10, -1.05847e-10, -1.060009e-10, -1.06438e-10, -1.068319e-10, 
    -1.072614e-10, -1.073665e-10, -1.078683e-10, -1.074598e-10, -1.08134e-10, 
    -1.075609e-10, -1.085529e-10, -1.067704e-10, -1.07544e-10, -1.061424e-10, 
    -1.062934e-10, -1.065665e-10, -1.071929e-10, -1.068547e-10, 
    -1.072502e-10, -1.063767e-10, -1.059236e-10, -1.058063e-10, 
    -1.055876e-10, -1.058113e-10, -1.057931e-10, -1.060072e-10, 
    -1.059384e-10, -1.064525e-10, -1.061764e-10, -1.069608e-10, 
    -1.072471e-10, -1.080555e-10, -1.085511e-10, -1.090555e-10, 
    -1.092782e-10, -1.09346e-10, -1.093744e-10 ;

 SMINN_TO_SOIL3N_S2 =
  -8.62019e-12, -8.658123e-12, -8.650748e-12, -8.681344e-12, -8.664371e-12, 
    -8.684406e-12, -8.62788e-12, -8.659629e-12, -8.639361e-12, -8.623604e-12, 
    -8.740719e-12, -8.682708e-12, -8.800973e-12, -8.763977e-12, 
    -8.856911e-12, -8.795216e-12, -8.869351e-12, -8.85513e-12, -8.897928e-12, 
    -8.885667e-12, -8.940411e-12, -8.903587e-12, -8.968787e-12, 
    -8.931616e-12, -8.937432e-12, -8.902373e-12, -8.694382e-12, 
    -8.733497e-12, -8.692064e-12, -8.697642e-12, -8.695139e-12, 
    -8.664722e-12, -8.649395e-12, -8.61729e-12, -8.623118e-12, -8.646698e-12, 
    -8.700151e-12, -8.682005e-12, -8.727734e-12, -8.726701e-12, 
    -8.777611e-12, -8.754657e-12, -8.840223e-12, -8.815904e-12, 
    -8.886179e-12, -8.868506e-12, -8.885349e-12, -8.880241e-12, 
    -8.885416e-12, -8.859496e-12, -8.870601e-12, -8.847792e-12, 
    -8.758956e-12, -8.785065e-12, -8.707196e-12, -8.660375e-12, 
    -8.629273e-12, -8.607203e-12, -8.610323e-12, -8.616271e-12, 
    -8.646836e-12, -8.675572e-12, -8.697471e-12, -8.71212e-12, -8.726552e-12, 
    -8.770244e-12, -8.793366e-12, -8.845141e-12, -8.835797e-12, 
    -8.851626e-12, -8.866748e-12, -8.892136e-12, -8.887957e-12, 
    -8.899143e-12, -8.851208e-12, -8.883066e-12, -8.830475e-12, 
    -8.844858e-12, -8.730481e-12, -8.6869e-12, -8.668379e-12, -8.652166e-12, 
    -8.612722e-12, -8.639961e-12, -8.629223e-12, -8.654769e-12, 
    -8.671001e-12, -8.662972e-12, -8.712519e-12, -8.693257e-12, 
    -8.794737e-12, -8.751027e-12, -8.864983e-12, -8.837714e-12, -8.87152e-12, 
    -8.85427e-12, -8.883827e-12, -8.857226e-12, -8.903305e-12, -8.91334e-12, 
    -8.906482e-12, -8.932821e-12, -8.85575e-12, -8.885349e-12, -8.662748e-12, 
    -8.664057e-12, -8.670157e-12, -8.643344e-12, -8.641704e-12, -8.61713e-12, 
    -8.638995e-12, -8.648306e-12, -8.671942e-12, -8.685923e-12, 
    -8.699212e-12, -8.728433e-12, -8.761067e-12, -8.806699e-12, 
    -8.839482e-12, -8.861457e-12, -8.847982e-12, -8.859879e-12, -8.84658e-12, 
    -8.840346e-12, -8.909581e-12, -8.870705e-12, -8.929034e-12, 
    -8.925805e-12, -8.899409e-12, -8.92617e-12, -8.664977e-12, -8.657442e-12, 
    -8.631282e-12, -8.651754e-12, -8.614454e-12, -8.635334e-12, 
    -8.647339e-12, -8.69366e-12, -8.703837e-12, -8.713274e-12, -8.731912e-12, 
    -8.755832e-12, -8.797792e-12, -8.8343e-12, -8.867627e-12, -8.865185e-12, 
    -8.866045e-12, -8.87349e-12, -8.855048e-12, -8.876518e-12, -8.880121e-12, 
    -8.870699e-12, -8.925373e-12, -8.909753e-12, -8.925737e-12, 
    -8.915567e-12, -8.659891e-12, -8.672569e-12, -8.665718e-12, 
    -8.678601e-12, -8.669525e-12, -8.709882e-12, -8.721981e-12, 
    -8.778597e-12, -8.755361e-12, -8.79234e-12, -8.759117e-12, -8.765004e-12, 
    -8.793548e-12, -8.760912e-12, -8.832287e-12, -8.783899e-12, 
    -8.873779e-12, -8.82546e-12, -8.876807e-12, -8.867483e-12, -8.882921e-12, 
    -8.896749e-12, -8.914143e-12, -8.94624e-12, -8.938808e-12, -8.965649e-12, 
    -8.691469e-12, -8.707914e-12, -8.706465e-12, -8.723675e-12, 
    -8.736401e-12, -8.763985e-12, -8.808228e-12, -8.79159e-12, -8.822132e-12, 
    -8.828264e-12, -8.781862e-12, -8.810353e-12, -8.718919e-12, 
    -8.733693e-12, -8.724896e-12, -8.692767e-12, -8.795425e-12, 
    -8.742741e-12, -8.840024e-12, -8.811484e-12, -8.894777e-12, 
    -8.853355e-12, -8.934716e-12, -8.9695e-12, -9.002232e-12, -9.040489e-12, 
    -8.716888e-12, -8.705714e-12, -8.725721e-12, -8.753401e-12, 
    -8.779082e-12, -8.813225e-12, -8.816718e-12, -8.823114e-12, 
    -8.839682e-12, -8.853612e-12, -8.825138e-12, -8.857104e-12, -8.73712e-12, 
    -8.799998e-12, -8.701491e-12, -8.731155e-12, -8.751769e-12, 
    -8.742725e-12, -8.789689e-12, -8.800757e-12, -8.845737e-12, 
    -8.822485e-12, -8.960915e-12, -8.89967e-12, -9.069615e-12, -9.022123e-12, 
    -8.70181e-12, -8.716849e-12, -8.769189e-12, -8.744286e-12, -8.815504e-12, 
    -8.833034e-12, -8.847284e-12, -8.865501e-12, -8.867468e-12, 
    -8.878261e-12, -8.860574e-12, -8.877562e-12, -8.813297e-12, 
    -8.842016e-12, -8.763206e-12, -8.782388e-12, -8.773563e-12, 
    -8.763885e-12, -8.793758e-12, -8.825586e-12, -8.826265e-12, 
    -8.836471e-12, -8.865232e-12, -8.815793e-12, -8.968822e-12, 
    -8.874317e-12, -8.733248e-12, -8.762217e-12, -8.766352e-12, 
    -8.755131e-12, -8.831277e-12, -8.803687e-12, -8.877998e-12, 
    -8.857914e-12, -8.890821e-12, -8.874469e-12, -8.872064e-12, 
    -8.851061e-12, -8.837986e-12, -8.804952e-12, -8.778073e-12, 
    -8.756758e-12, -8.761714e-12, -8.785129e-12, -8.827532e-12, 
    -8.867646e-12, -8.858859e-12, -8.88832e-12, -8.81034e-12, -8.843039e-12, 
    -8.830402e-12, -8.863354e-12, -8.791148e-12, -8.852639e-12, 
    -8.775431e-12, -8.782201e-12, -8.803139e-12, -8.845258e-12, 
    -8.854574e-12, -8.864525e-12, -8.858385e-12, -8.828609e-12, -8.82373e-12, 
    -8.80263e-12, -8.796804e-12, -8.780726e-12, -8.767416e-12, -8.779578e-12, 
    -8.79235e-12, -8.828621e-12, -8.861308e-12, -8.896946e-12, -8.905666e-12, 
    -8.947308e-12, -8.913412e-12, -8.969349e-12, -8.921794e-12, 
    -9.004113e-12, -8.8562e-12, -8.920393e-12, -8.804091e-12, -8.816621e-12, 
    -8.839283e-12, -8.891261e-12, -8.863198e-12, -8.896017e-12, 
    -8.823539e-12, -8.785937e-12, -8.776206e-12, -8.758055e-12, 
    -8.776622e-12, -8.775112e-12, -8.792878e-12, -8.787169e-12, 
    -8.829825e-12, -8.806912e-12, -8.872003e-12, -8.895757e-12, 
    -8.962837e-12, -9.003959e-12, -9.045817e-12, -9.064297e-12, 
    -9.069922e-12, -9.072273e-12 ;

 SMIN_NH4 =
  0.0004618175, 0.0004637462, 0.0004633711, 0.0004649268, 0.0004640637, 
    0.0004650823, 0.0004622081, 0.0004638225, 0.0004627918, 0.0004619905, 
    0.0004679451, 0.0004649957, 0.0004710071, 0.0004691266, 0.0004738494, 
    0.0004707145, 0.0004744813, 0.0004737586, 0.0004759328, 0.0004753099, 
    0.000478091, 0.0004762202, 0.000479532, 0.000477644, 0.0004779394, 
    0.0004761582, 0.0004655895, 0.0004675784, 0.0004654716, 0.0004657552, 
    0.0004656278, 0.0004640814, 0.0004633022, 0.0004616693, 0.0004619657, 
    0.0004631648, 0.0004658824, 0.0004649597, 0.0004672842, 0.0004672317, 
    0.0004698193, 0.0004686527, 0.0004730011, 0.0004717651, 0.0004753358, 
    0.0004744379, 0.0004752936, 0.000475034, 0.0004752968, 0.0004739799, 
    0.0004745441, 0.0004733852, 0.0004688719, 0.0004701988, 0.0004662407, 
    0.0004638605, 0.0004622788, 0.0004611565, 0.000461315, 0.0004616175, 
    0.0004631717, 0.0004646325, 0.0004657458, 0.0004664904, 0.000467224, 
    0.0004694453, 0.0004706201, 0.000473251, 0.000472776, 0.0004735803, 
    0.0004743485, 0.0004756383, 0.0004754259, 0.0004759941, 0.0004735587, 
    0.0004751774, 0.000472505, 0.000473236, 0.0004674249, 0.0004652088, 
    0.0004642674, 0.0004634428, 0.000461437, 0.0004628222, 0.0004622761, 
    0.0004635748, 0.0004644001, 0.0004639918, 0.0004665107, 0.0004655314, 
    0.0004706897, 0.0004684681, 0.000474259, 0.0004728733, 0.0004745908, 
    0.0004737144, 0.0004752161, 0.0004738645, 0.0004762055, 0.0004767153, 
    0.0004763668, 0.0004777047, 0.0004737892, 0.0004752931, 0.0004639807, 
    0.0004640473, 0.0004643573, 0.0004629941, 0.0004629106, 0.0004616609, 
    0.0004627727, 0.0004632462, 0.0004644477, 0.0004651585, 0.0004658341, 
    0.0004673195, 0.0004689783, 0.0004712974, 0.0004729631, 0.0004740795, 
    0.0004733948, 0.0004739992, 0.0004733235, 0.0004730066, 0.0004765242, 
    0.0004745492, 0.0004775121, 0.0004773482, 0.0004760073, 0.0004773665, 
    0.0004640939, 0.0004637107, 0.0004623806, 0.0004634215, 0.0004615247, 
    0.0004625865, 0.000463197, 0.000465552, 0.0004660691, 0.0004665489, 
    0.0004674962, 0.000468712, 0.0004708446, 0.0004726997, 0.0004743929, 
    0.0004742687, 0.0004743124, 0.0004746907, 0.0004737536, 0.0004748444, 
    0.0004750274, 0.0004745487, 0.000477326, 0.0004765326, 0.0004773445, 
    0.0004768277, 0.0004638352, 0.0004644797, 0.0004641313, 0.0004647864, 
    0.0004643248, 0.0004663767, 0.0004669917, 0.0004698693, 0.0004686881, 
    0.0004705676, 0.0004688788, 0.0004691781, 0.0004706291, 0.0004689699, 
    0.0004725974, 0.0004701384, 0.0004747053, 0.0004722504, 0.000474859, 
    0.0004743851, 0.0004751694, 0.000475872, 0.0004767555, 0.000478386, 
    0.0004780083, 0.0004793716, 0.0004654406, 0.0004662766, 0.0004662028, 
    0.0004670775, 0.0004677244, 0.0004691264, 0.0004713749, 0.0004705293, 
    0.0004720813, 0.0004723929, 0.0004700347, 0.0004714827, 0.0004668354, 
    0.0004675864, 0.0004671391, 0.0004655058, 0.0004707239, 0.0004680462, 
    0.00047299, 0.0004715396, 0.0004757717, 0.0004736673, 0.0004778004, 
    0.0004795674, 0.0004812293, 0.0004831721, 0.0004667326, 0.0004661645, 
    0.0004671814, 0.0004685886, 0.0004698936, 0.0004716288, 0.0004718061, 
    0.0004721311, 0.0004729729, 0.0004736807, 0.0004722339, 0.000473858, 
    0.0004677609, 0.0004709562, 0.0004659491, 0.0004674573, 0.0004685048, 
    0.0004680451, 0.0004704319, 0.0004709943, 0.00047328, 0.0004720984, 
    0.0004791313, 0.0004760202, 0.0004846506, 0.0004822394, 0.000465966, 
    0.0004667304, 0.0004693909, 0.000468125, 0.0004717444, 0.0004726352, 
    0.0004733591, 0.0004742848, 0.0004743845, 0.000474933, 0.0004740342, 
    0.0004748973, 0.0004716319, 0.0004730912, 0.000469086, 0.0004700609, 
    0.0004696123, 0.0004691203, 0.0004706385, 0.0004722561, 0.0004722904, 
    0.000472809, 0.000474271, 0.000471758, 0.000479533, 0.0004747322, 
    0.0004675639, 0.0004690365, 0.0004692464, 0.0004686761, 0.0004725458, 
    0.0004711438, 0.0004749196, 0.000473899, 0.0004755708, 0.0004747401, 
    0.0004746178, 0.0004735507, 0.0004728863, 0.0004712077, 0.0004698415, 
    0.0004687581, 0.0004690099, 0.0004702, 0.0004723548, 0.000474393, 
    0.0004739465, 0.0004754431, 0.0004714808, 0.0004731425, 0.0004725003, 
    0.0004741745, 0.0004705066, 0.0004736319, 0.0004697077, 0.0004700517, 
    0.0004711158, 0.0004732563, 0.0004737292, 0.0004742349, 0.0004739227, 
    0.0004724099, 0.0004721619, 0.0004710895, 0.0004707935, 0.0004699763, 
    0.0004692996, 0.0004699178, 0.0004705669, 0.00047241, 0.0004740709, 
    0.0004758813, 0.0004763243, 0.0004784398, 0.0004767179, 0.0004795596, 
    0.0004771441, 0.0004813247, 0.0004738124, 0.0004770737, 0.0004711641, 
    0.0004718007, 0.0004729525, 0.0004755933, 0.0004741673, 0.0004758348, 
    0.0004721521, 0.0004702413, 0.0004697465, 0.0004688239, 0.0004697675, 
    0.0004696907, 0.0004705936, 0.0004703033, 0.0004724711, 0.0004713066, 
    0.0004746141, 0.0004758209, 0.0004792282, 0.0004813166, 0.0004834418, 
    0.00048438, 0.0004846655, 0.0004847849 ;

 SMIN_NH4_vr =
  0.00302471, 0.003029867, 0.003028858, 0.003033014, 0.003030704, 
    0.003033421, 0.003025739, 0.003030051, 0.003027294, 0.003025146, 
    0.003041045, 0.003033175, 0.003049191, 0.003044181, 0.003056736, 
    0.003048406, 0.00305841, 0.003056486, 0.003062254, 0.003060597, 
    0.003067966, 0.003063007, 0.003071774, 0.003066776, 0.003067555, 
    0.003062829, 0.00303478, 0.00304009, 0.003034459, 0.003035217, 
    0.003034873, 0.00303074, 0.003028658, 0.003024285, 0.003025074, 
    0.003028281, 0.003035535, 0.003033067, 0.003039265, 0.003039125, 
    0.003046013, 0.003042907, 0.003054471, 0.003051181, 0.003060662, 
    0.003058275, 0.003060544, 0.003059851, 0.003060544, 0.003057051, 
    0.003058542, 0.003055465, 0.003043526, 0.003047054, 0.003036506, 
    0.003030149, 0.003025916, 0.003022914, 0.003023332, 0.003024142, 
    0.003028294, 0.003032191, 0.003035162, 0.003037144, 0.003039096, 
    0.003045018, 0.00304814, 0.003055128, 0.003053864, 0.003055997, 
    0.003058034, 0.003061452, 0.003060887, 0.00306239, 0.003055923, 
    0.003060221, 0.003053118, 0.003055061, 0.003039666, 0.003033745, 
    0.003031233, 0.003029023, 0.003023656, 0.003027362, 0.003025898, 
    0.003029364, 0.003031567, 0.003030472, 0.003037194, 0.003034577, 
    0.00304832, 0.003042405, 0.003057801, 0.003054116, 0.003058673, 
    0.003056347, 0.003060326, 0.003056739, 0.003062944, 0.003064297, 
    0.003063367, 0.003066912, 0.003056521, 0.003060514, 0.00303046, 
    0.003030639, 0.003031463, 0.003027817, 0.003027592, 0.003024245, 
    0.003027214, 0.003028481, 0.003031686, 0.00303358, 0.003035379, 
    0.003039342, 0.003043759, 0.003049926, 0.003054351, 0.003057311, 
    0.003055492, 0.003057092, 0.003055297, 0.00305445, 0.003063782, 
    0.003058544, 0.003066393, 0.003065959, 0.003062402, 0.003065999, 
    0.003030757, 0.003029728, 0.003026173, 0.00302895, 0.003023874, 
    0.003026715, 0.003028344, 0.003034629, 0.003036004, 0.003037285, 
    0.003039807, 0.003043042, 0.003048718, 0.003053645, 0.00305814, 
    0.003057806, 0.00305792, 0.00305892, 0.003056431, 0.003059322, 
    0.003059804, 0.003058534, 0.003065892, 0.00306379, 0.003065938, 
    0.003064564, 0.003030058, 0.003031775, 0.00303084, 0.003032591, 
    0.003031352, 0.00303683, 0.003038467, 0.003046129, 0.003042978, 
    0.003047983, 0.00304348, 0.003044278, 0.003048139, 0.003043715, 
    0.003053366, 0.003046822, 0.003058956, 0.003052434, 0.003059358, 
    0.003058095, 0.003060172, 0.003062037, 0.003064372, 0.003068693, 
    0.003067686, 0.003071295, 0.003034337, 0.003036564, 0.003036365, 
    0.003038693, 0.003040414, 0.00304415, 0.00305013, 0.003047875, 
    0.003051999, 0.003052828, 0.003046549, 0.003050403, 0.003038024, 
    0.003040022, 0.003038827, 0.003034466, 0.00304837, 0.003041236, 
    0.003054387, 0.003050528, 0.003061762, 0.003056179, 0.003067133, 
    0.003071813, 0.003076201, 0.00308133, 0.003037776, 0.003036256, 
    0.003038964, 0.003042717, 0.003046184, 0.003050801, 0.003051268, 
    0.003052128, 0.00305436, 0.003056241, 0.003052395, 0.003056703, 
    0.003040486, 0.003048987, 0.003035643, 0.003039667, 0.003042451, 
    0.003041227, 0.003047577, 0.003049069, 0.003055142, 0.003052002, 
    0.003070651, 0.00306241, 0.003085223, 0.003078862, 0.003035723, 
    0.003037757, 0.003044844, 0.003041473, 0.003051099, 0.003053468, 
    0.003055384, 0.003057844, 0.003058101, 0.003059558, 0.003057165, 
    0.003059457, 0.003050777, 0.003054656, 0.003043998, 0.00304659, 
    0.003045394, 0.00304408, 0.003048117, 0.003052421, 0.003052506, 
    0.003053881, 0.003057767, 0.003051081, 0.003071706, 0.00305898, 
    0.003039977, 0.003043897, 0.003044451, 0.003042932, 0.003053222, 
    0.003049495, 0.003059522, 0.003056808, 0.003061241, 0.003059037, 
    0.003058706, 0.003055874, 0.003054103, 0.003049642, 0.003046, 
    0.003043115, 0.003043779, 0.003046949, 0.003052674, 0.003058088, 
    0.003056899, 0.003060865, 0.003050338, 0.003054756, 0.003053043, 
    0.00305749, 0.003047803, 0.003056116, 0.003045673, 0.003046584, 
    0.003049412, 0.003055104, 0.003056351, 0.003057695, 0.003056859, 
    0.003052842, 0.003052179, 0.003049322, 0.003048531, 0.003046357, 
    0.003044549, 0.003046196, 0.003047917, 0.003052818, 0.003057227, 
    0.003062025, 0.003063198, 0.003068802, 0.003064238, 0.003071762, 
    0.003065365, 0.003076421, 0.003056585, 0.003065236, 0.003049541, 
    0.003051229, 0.00305429, 0.003061296, 0.003057507, 0.003061933, 
    0.00305215, 0.003047065, 0.003045743, 0.003043287, 0.003045792, 
    0.003045589, 0.003047988, 0.003047211, 0.003052972, 0.003049877, 
    0.003058658, 0.003061861, 0.003070883, 0.003076401, 0.00308201, 
    0.003084481, 0.003085232, 0.003085543,
  0.00181022, 0.001816974, 0.001815662, 0.001821105, 0.001818086, 0.00182165, 
    0.00181159, 0.001817243, 0.001813634, 0.001810828, 0.001831657, 
    0.001821348, 0.001842343, 0.001835782, 0.001852247, 0.001841323, 
    0.001854447, 0.001851931, 0.001859498, 0.001857331, 0.001867001, 
    0.001860497, 0.001872005, 0.001865448, 0.001866474, 0.001860283, 
    0.001823423, 0.001830375, 0.001823011, 0.001824003, 0.001823558, 
    0.001818148, 0.001815422, 0.001809703, 0.001810741, 0.001814941, 
    0.001824449, 0.001821222, 0.001829349, 0.001829165, 0.0018382, 
    0.001834128, 0.001849293, 0.001844987, 0.001857421, 0.001854297, 
    0.001857275, 0.001856372, 0.001857287, 0.001852703, 0.001854668, 
    0.001850633, 0.001834891, 0.001839522, 0.001825701, 0.001817376, 
    0.001811838, 0.001807906, 0.001808462, 0.001809522, 0.001814965, 
    0.001820078, 0.001823972, 0.001826575, 0.001829139, 0.001836895, 
    0.001840994, 0.001850164, 0.001848509, 0.001851311, 0.001853986, 
    0.001858474, 0.001857736, 0.001859713, 0.001851237, 0.001856872, 
    0.001847567, 0.001850113, 0.001829839, 0.001822093, 0.0018188, 
    0.001815914, 0.00180889, 0.001813742, 0.001811829, 0.001816377, 
    0.001819265, 0.001817837, 0.001826646, 0.001823223, 0.001841237, 
    0.001833485, 0.001853674, 0.001848849, 0.00185483, 0.001851778, 
    0.001857006, 0.001852301, 0.001860448, 0.001862221, 0.001861009, 
    0.00186566, 0.001852041, 0.001857275, 0.001817797, 0.00181803, 
    0.001819115, 0.001814344, 0.001814052, 0.001809675, 0.001813569, 
    0.001815227, 0.001819432, 0.001821919, 0.001824282, 0.001829473, 
    0.001835266, 0.001843357, 0.001849162, 0.00185305, 0.001850666, 
    0.001852771, 0.001850418, 0.001849315, 0.001861557, 0.001854686, 
    0.001864991, 0.001864421, 0.00185976, 0.001864486, 0.001818193, 
    0.001816852, 0.001812196, 0.00181584, 0.001809198, 0.001812917, 
    0.001815055, 0.001823295, 0.001825103, 0.00182678, 0.001830091, 
    0.001834337, 0.001841778, 0.001848245, 0.001854141, 0.001853709, 
    0.001853861, 0.001855178, 0.001851916, 0.001855714, 0.001856351, 
    0.001854685, 0.001864345, 0.001861587, 0.001864409, 0.001862613, 
    0.001817288, 0.001819544, 0.001818325, 0.001820617, 0.001819003, 
    0.001826178, 0.001828328, 0.001838376, 0.001834253, 0.001840812, 
    0.00183492, 0.001835964, 0.001841028, 0.001835238, 0.001847889, 
    0.001839316, 0.001855229, 0.001846681, 0.001855765, 0.001854116, 
    0.001856845, 0.00185929, 0.001862362, 0.001868028, 0.001866717, 
    0.001871451, 0.001822905, 0.001825828, 0.00182557, 0.001828628, 
    0.001830888, 0.001835783, 0.001843627, 0.001840679, 0.00184609, 
    0.001847176, 0.001838954, 0.001844004, 0.001827783, 0.001830408, 
    0.001828845, 0.001823136, 0.001841359, 0.001832014, 0.001849258, 
    0.001844204, 0.001858941, 0.001851617, 0.001865995, 0.001872131, 
    0.001877898, 0.001884633, 0.001827422, 0.001825437, 0.001828991, 
    0.001833906, 0.001838461, 0.001844513, 0.001845131, 0.001846264, 
    0.001849197, 0.001851662, 0.001846623, 0.00185228, 0.001831018, 
    0.001842169, 0.001824687, 0.001829957, 0.001833616, 0.001832011, 
    0.001840341, 0.001842303, 0.001850269, 0.001846152, 0.001870618, 
    0.001859807, 0.001889753, 0.001881401, 0.001824743, 0.001827415, 
    0.001836707, 0.001832288, 0.001844916, 0.00184802, 0.001850542, 
    0.001853766, 0.001854113, 0.001856022, 0.001852894, 0.001855898, 
    0.001844525, 0.00184961, 0.001835645, 0.001839047, 0.001837482, 
    0.001835765, 0.001841063, 0.001846702, 0.001846822, 0.001848629, 
    0.001853721, 0.001844967, 0.001872014, 0.001855327, 0.001830328, 
    0.001835471, 0.001836203, 0.001834212, 0.001847709, 0.001842823, 
    0.001855975, 0.001852423, 0.001858242, 0.001855351, 0.001854926, 
    0.001851211, 0.001848897, 0.001843047, 0.001838282, 0.001834501, 
    0.00183538, 0.001839533, 0.001847047, 0.001854145, 0.001852591, 
    0.0018578, 0.001844001, 0.001849792, 0.001847555, 0.001853386, 0.0018406, 
    0.001851493, 0.001837813, 0.001839014, 0.001842725, 0.001850185, 
    0.001851832, 0.001853593, 0.001852506, 0.001847237, 0.001846373, 
    0.001842635, 0.001841603, 0.001838752, 0.001836392, 0.001838549, 
    0.001840814, 0.001847239, 0.001853024, 0.001859325, 0.001860865, 
    0.001868218, 0.001862235, 0.001872107, 0.001863717, 0.001878231, 
    0.001852122, 0.001863468, 0.001842894, 0.001845114, 0.001849127, 
    0.001858321, 0.001853358, 0.001859161, 0.001846339, 0.001839677, 
    0.001837951, 0.001834731, 0.001838024, 0.001837757, 0.001840907, 
    0.001839894, 0.001847452, 0.001843394, 0.001854916, 0.001859115, 
    0.001870956, 0.001878203, 0.001885568, 0.001888818, 0.001889806, 
    0.001890219,
  0.001646094, 0.001653298, 0.001651898, 0.001657706, 0.001654484, 
    0.001658287, 0.001647554, 0.001653584, 0.001649735, 0.001646742, 
    0.001668967, 0.001657964, 0.001680378, 0.001673372, 0.00169096, 
    0.001679289, 0.001693311, 0.001690623, 0.00169871, 0.001696394, 
    0.001706732, 0.001699779, 0.001712085, 0.001705072, 0.00170617, 
    0.00169955, 0.001660179, 0.001667598, 0.001659739, 0.001660798, 
    0.001660323, 0.001654551, 0.001651641, 0.001645542, 0.00164665, 
    0.001651129, 0.001661274, 0.001657831, 0.001666504, 0.001666308, 
    0.001675955, 0.001671606, 0.001687804, 0.001683203, 0.001696491, 
    0.001693151, 0.001696334, 0.001695369, 0.001696347, 0.001691448, 
    0.001693547, 0.001689235, 0.001672421, 0.001677366, 0.00166261, 
    0.001653726, 0.001647819, 0.001643626, 0.001644219, 0.001645349, 
    0.001651155, 0.00165661, 0.001660765, 0.001663543, 0.00166628, 
    0.00167456, 0.001678938, 0.001688735, 0.001686967, 0.001689961, 
    0.001692819, 0.001697617, 0.001696827, 0.00169894, 0.001689881, 
    0.001695903, 0.00168596, 0.001688681, 0.001667026, 0.00165876, 
    0.001655246, 0.001652167, 0.001644675, 0.001649849, 0.00164781, 
    0.001652661, 0.001655742, 0.001654218, 0.001663619, 0.001659966, 
    0.001679198, 0.001670919, 0.001692486, 0.001687329, 0.001693721, 
    0.00169046, 0.001696047, 0.001691019, 0.001699726, 0.001701621, 
    0.001700326, 0.001705299, 0.00169074, 0.001696334, 0.001654176, 
    0.001654424, 0.001655582, 0.001650492, 0.00165018, 0.001645512, 
    0.001649666, 0.001651434, 0.001655921, 0.001658574, 0.001661095, 
    0.001666637, 0.001672821, 0.001681462, 0.001687664, 0.001691819, 
    0.001689271, 0.00169152, 0.001689006, 0.001687827, 0.001700912, 
    0.001693567, 0.001704584, 0.001703975, 0.00169899, 0.001704043, 
    0.001654599, 0.001653168, 0.001648201, 0.001652089, 0.001645004, 
    0.00164897, 0.001651251, 0.001660043, 0.001661972, 0.001663762, 
    0.001667296, 0.001671829, 0.001679776, 0.001686684, 0.001692985, 
    0.001692524, 0.001692686, 0.001694093, 0.001690607, 0.001694666, 
    0.001695347, 0.001693566, 0.001703893, 0.001700944, 0.001703962, 
    0.001702041, 0.001653633, 0.00165604, 0.00165474, 0.001657185, 
    0.001655462, 0.00166312, 0.001665414, 0.001676142, 0.00167174, 
    0.001678744, 0.001672452, 0.001673567, 0.001678973, 0.001672792, 
    0.001686304, 0.001677146, 0.001694148, 0.001685012, 0.00169472, 
    0.001692958, 0.001695875, 0.001698488, 0.001701773, 0.001707832, 
    0.001706429, 0.001711493, 0.001659626, 0.001662746, 0.001662471, 
    0.001665734, 0.001668147, 0.001673374, 0.001681751, 0.001678601, 
    0.001684382, 0.001685542, 0.00167676, 0.001682153, 0.001664833, 
    0.001667634, 0.001665966, 0.001659873, 0.001679328, 0.001669349, 
    0.001687767, 0.001682367, 0.001698115, 0.001690288, 0.001705657, 
    0.00171222, 0.001718389, 0.001725596, 0.001664448, 0.001662328, 
    0.001666122, 0.001671369, 0.001676233, 0.001682697, 0.001683357, 
    0.001684568, 0.001687702, 0.001690336, 0.001684951, 0.001690996, 
    0.001668285, 0.001680193, 0.001661528, 0.001667153, 0.00167106, 
    0.001669346, 0.001678241, 0.001680337, 0.001688847, 0.001684448, 
    0.001710601, 0.00169904, 0.001731078, 0.001722138, 0.001661588, 
    0.00166444, 0.00167436, 0.001669641, 0.001683128, 0.001686444, 
    0.001689139, 0.001692584, 0.001692955, 0.001694995, 0.001691652, 
    0.001694863, 0.00168271, 0.001688143, 0.001673226, 0.001676859, 
    0.001675188, 0.001673354, 0.001679012, 0.001685036, 0.001685164, 
    0.001687094, 0.001692535, 0.001683182, 0.001712093, 0.001694251, 
    0.001667549, 0.001673039, 0.001673822, 0.001671696, 0.001686112, 
    0.001680891, 0.001694945, 0.001691149, 0.001697368, 0.001694278, 
    0.001693824, 0.001689853, 0.001687381, 0.001681131, 0.001676042, 
    0.001672004, 0.001672943, 0.001677378, 0.001685404, 0.001692989, 
    0.001691328, 0.001696895, 0.00168215, 0.001688337, 0.001685946, 
    0.001692177, 0.001678518, 0.001690154, 0.001675542, 0.001676823, 
    0.001680788, 0.001688757, 0.001690518, 0.001692399, 0.001691238, 
    0.001685607, 0.001684684, 0.001680691, 0.001679589, 0.001676544, 
    0.001674023, 0.001676327, 0.001678745, 0.001685609, 0.001691791, 
    0.001698525, 0.001700172, 0.001708034, 0.001701636, 0.001712193, 
    0.00170322, 0.001718745, 0.001690826, 0.001702954, 0.001680968, 
    0.001683339, 0.001687627, 0.001697452, 0.001692148, 0.00169835, 
    0.001684648, 0.001677532, 0.001675688, 0.00167225, 0.001675767, 
    0.001675481, 0.001678845, 0.001677764, 0.001685837, 0.001681502, 
    0.001693812, 0.001698301, 0.001710963, 0.001718715, 0.001726599, 
    0.001730077, 0.001731135, 0.001731578,
  0.001514893, 0.001522024, 0.001520637, 0.001526388, 0.001523198, 
    0.001526964, 0.001516338, 0.001522307, 0.001518497, 0.001515534, 
    0.001537545, 0.001526645, 0.00154886, 0.001541913, 0.001559361, 
    0.00154778, 0.001561695, 0.001559026, 0.001567057, 0.001564757, 
    0.001575027, 0.001568119, 0.001580348, 0.001573377, 0.001574468, 
    0.001567891, 0.001528838, 0.001536189, 0.001528403, 0.001529451, 
    0.00152898, 0.001523264, 0.001520383, 0.001514347, 0.001515443, 
    0.001519876, 0.001529922, 0.001526512, 0.001535104, 0.00153491, 
    0.001544473, 0.001540162, 0.001556228, 0.001551663, 0.001564853, 
    0.001561536, 0.001564697, 0.001563739, 0.001564709, 0.001559846, 
    0.00156193, 0.001557649, 0.001540969, 0.001545873, 0.001531246, 
    0.001522448, 0.0015166, 0.001512451, 0.001513037, 0.001514156, 
    0.001519902, 0.001525303, 0.001529418, 0.001532171, 0.001534882, 
    0.00154309, 0.001547432, 0.001557152, 0.001555397, 0.001558369, 
    0.001561206, 0.00156597, 0.001565186, 0.001567285, 0.00155829, 
    0.001564269, 0.001554398, 0.001557098, 0.001535622, 0.001527432, 
    0.001523952, 0.001520904, 0.001513488, 0.00151861, 0.001516591, 
    0.001521393, 0.001524444, 0.001522935, 0.001532246, 0.001528627, 
    0.001547689, 0.00153948, 0.001560875, 0.001555757, 0.001562102, 
    0.001558865, 0.001564412, 0.001559419, 0.001568066, 0.001569949, 
    0.001568662, 0.001573603, 0.001559143, 0.001564697, 0.001522893, 
    0.001523139, 0.001524285, 0.001519246, 0.001518937, 0.001514317, 
    0.001518428, 0.001520178, 0.001524621, 0.001527248, 0.001529746, 
    0.001535236, 0.001541366, 0.001549935, 0.001556089, 0.001560214, 
    0.001557685, 0.001559917, 0.001557421, 0.001556251, 0.001569243, 
    0.001561949, 0.001572892, 0.001572287, 0.001567335, 0.001572355, 
    0.001523312, 0.001521895, 0.001516978, 0.001520826, 0.001513814, 
    0.00151774, 0.001519997, 0.001528703, 0.001530615, 0.001532388, 
    0.001535889, 0.001540383, 0.001548263, 0.001555117, 0.001561371, 
    0.001560913, 0.001561075, 0.001562472, 0.001559011, 0.00156304, 
    0.001563716, 0.001561948, 0.001572206, 0.001569276, 0.001572274, 
    0.001570366, 0.001522356, 0.001524739, 0.001523451, 0.001525873, 
    0.001524167, 0.001531751, 0.001534024, 0.001544659, 0.001540294, 
    0.001547239, 0.001541, 0.001542106, 0.001547467, 0.001541337, 
    0.001554739, 0.001545654, 0.001562526, 0.001553458, 0.001563094, 
    0.001561344, 0.001564241, 0.001566836, 0.001570099, 0.00157612, 
    0.001574725, 0.001579759, 0.001528291, 0.001531381, 0.001531108, 
    0.001534342, 0.001536733, 0.001541914, 0.001550222, 0.001547098, 
    0.001552832, 0.001553983, 0.001545271, 0.001550621, 0.001533449, 
    0.001536224, 0.001534571, 0.001528535, 0.001547819, 0.001537924, 
    0.001556191, 0.001550833, 0.001566466, 0.001558693, 0.001573958, 
    0.001580482, 0.001586618, 0.001593788, 0.001533067, 0.001530967, 
    0.001534726, 0.001539927, 0.001544749, 0.00155116, 0.001551816, 
    0.001553017, 0.001556127, 0.001558741, 0.001553397, 0.001559397, 
    0.001536869, 0.001548677, 0.001530174, 0.001535748, 0.00153962, 
    0.001537921, 0.001546741, 0.001548819, 0.001557264, 0.001552898, 
    0.001578872, 0.001567384, 0.001599245, 0.001590346, 0.001530234, 
    0.001533059, 0.001542892, 0.001538214, 0.001551588, 0.001554879, 
    0.001557554, 0.001560973, 0.001561342, 0.001563367, 0.001560048, 
    0.001563236, 0.001551174, 0.001556565, 0.001541768, 0.00154537, 
    0.001543713, 0.001541895, 0.001547505, 0.001553481, 0.001553608, 
    0.001555524, 0.001560924, 0.001551642, 0.001580356, 0.001562629, 
    0.00153614, 0.001541582, 0.001542359, 0.001540251, 0.001554549, 
    0.001549369, 0.001563318, 0.001559549, 0.001565724, 0.001562655, 
    0.001562204, 0.001558263, 0.001555808, 0.001549607, 0.00154456, 
    0.001540557, 0.001541487, 0.001545885, 0.001553847, 0.001561375, 
    0.001559726, 0.001565254, 0.001550618, 0.001556757, 0.001554385, 
    0.00156057, 0.001547015, 0.00155856, 0.001544063, 0.001545335, 
    0.001549267, 0.001557174, 0.001558922, 0.001560789, 0.001559637, 
    0.001554048, 0.001553132, 0.001549171, 0.001548077, 0.001545058, 
    0.001542558, 0.001544842, 0.001547241, 0.00155405, 0.001560186, 
    0.001566873, 0.001568509, 0.001576321, 0.001569963, 0.001580455, 
    0.001571536, 0.001586972, 0.001559228, 0.001571273, 0.001549445, 
    0.001551797, 0.001556052, 0.001565807, 0.001560541, 0.001566699, 
    0.001553096, 0.001546037, 0.001544209, 0.0015408, 0.001544287, 
    0.001544003, 0.00154734, 0.001546268, 0.001554277, 0.001549975, 
    0.001562193, 0.00156665, 0.001579232, 0.001586942, 0.001594786, 
    0.001598249, 0.001599302, 0.001599743,
  0.0013795, 0.001385892, 0.001384649, 0.001389807, 0.001386945, 0.001390323, 
    0.001380795, 0.001386146, 0.00138273, 0.001380075, 0.001399825, 
    0.001390037, 0.001409999, 0.00140375, 0.001419454, 0.001409026, 
    0.001421557, 0.001419152, 0.001426391, 0.001424317, 0.001433584, 
    0.001427349, 0.00143839, 0.001432094, 0.001433079, 0.001427144, 
    0.001392005, 0.001398606, 0.001391615, 0.001392556, 0.001392133, 
    0.001387005, 0.001384421, 0.001379011, 0.001379993, 0.001383967, 
    0.001392979, 0.001389918, 0.001397632, 0.001397458, 0.001406052, 
    0.001402176, 0.001416632, 0.001412521, 0.001424404, 0.001421414, 
    0.001424263, 0.001423399, 0.001424274, 0.00141989, 0.001421768, 
    0.001417911, 0.001402902, 0.001407311, 0.001394167, 0.001386272, 
    0.00138103, 0.001377312, 0.001377838, 0.00137884, 0.00138399, 
    0.001388833, 0.001392526, 0.001394997, 0.001397433, 0.001404809, 
    0.001408714, 0.001417463, 0.001415883, 0.00141856, 0.001421117, 
    0.001425412, 0.001424704, 0.001426597, 0.001418489, 0.001423877, 
    0.001414983, 0.001417415, 0.001398097, 0.001390744, 0.001387622, 
    0.001384888, 0.001378242, 0.001382831, 0.001381022, 0.001385326, 
    0.001388063, 0.001386709, 0.001395065, 0.001391816, 0.001408945, 
    0.001401564, 0.001420818, 0.001416207, 0.001421924, 0.001419006, 
    0.001424006, 0.001419506, 0.001427302, 0.001429, 0.001427839, 
    0.001432298, 0.001419257, 0.001424263, 0.001386671, 0.001386892, 
    0.00138792, 0.001383401, 0.001383125, 0.001378985, 0.001382668, 
    0.001384238, 0.001388221, 0.001390579, 0.00139282, 0.00139775, 
    0.001403259, 0.001410966, 0.001416506, 0.001420222, 0.001417943, 
    0.001419955, 0.001417706, 0.001416652, 0.001428364, 0.001421786, 
    0.001431657, 0.00143111, 0.001426642, 0.001431172, 0.001387047, 
    0.001385777, 0.001381369, 0.001384818, 0.001378534, 0.001382051, 
    0.001384075, 0.001391884, 0.0013936, 0.001395192, 0.001398337, 
    0.001402374, 0.001409461, 0.00141563, 0.001421265, 0.001420852, 
    0.001420998, 0.001422257, 0.001419138, 0.001422769, 0.001423379, 
    0.001421785, 0.001431037, 0.001428393, 0.001431098, 0.001429377, 
    0.00138619, 0.001388327, 0.001387172, 0.001389344, 0.001387814, 
    0.00139462, 0.001396662, 0.001406219, 0.001402295, 0.00140854, 
    0.001402929, 0.001403923, 0.001408745, 0.001403232, 0.001415291, 
    0.001407115, 0.001422306, 0.001414137, 0.001422818, 0.001421241, 
    0.001423852, 0.001426192, 0.001429136, 0.001434571, 0.001433312, 
    0.001437858, 0.001391514, 0.001394288, 0.001394044, 0.001396947, 
    0.001399095, 0.001403751, 0.001411224, 0.001408413, 0.001413573, 
    0.00141461, 0.00140677, 0.001411583, 0.001396145, 0.001398638, 
    0.001397153, 0.001391733, 0.001409061, 0.001400165, 0.001416598, 
    0.001411774, 0.001425858, 0.001418852, 0.001432619, 0.001438511, 
    0.001444058, 0.001450546, 0.001395802, 0.001393917, 0.001397292, 
    0.001401965, 0.0014063, 0.001412068, 0.001412658, 0.00141374, 0.00141654, 
    0.001418895, 0.001414082, 0.001419486, 0.001399217, 0.001409834, 
    0.001393205, 0.00139821, 0.001401689, 0.001400162, 0.001408092, 
    0.001409962, 0.001417564, 0.001413633, 0.001437057, 0.001426687, 
    0.001455488, 0.001447431, 0.001393258, 0.001395795, 0.00140463, 
    0.001400425, 0.001412453, 0.001415416, 0.001417825, 0.001420906, 
    0.001421238, 0.001423064, 0.001420072, 0.001422946, 0.001412081, 
    0.001416935, 0.001403619, 0.001406859, 0.001405368, 0.001403734, 
    0.001408779, 0.001414158, 0.001414272, 0.001415997, 0.001420862, 
    0.001412502, 0.001438398, 0.001422399, 0.001398562, 0.001403453, 
    0.001404151, 0.001402256, 0.001415119, 0.001410457, 0.00142302, 
    0.001419623, 0.001425189, 0.001422423, 0.001422016, 0.001418464, 
    0.001416253, 0.001410671, 0.00140613, 0.001402531, 0.001403367, 
    0.001407322, 0.001414487, 0.001421269, 0.001419783, 0.001424766, 
    0.001411581, 0.001417108, 0.001414971, 0.001420543, 0.001408338, 
    0.001418732, 0.001405684, 0.001406827, 0.001410364, 0.001417483, 
    0.001419058, 0.001420741, 0.001419702, 0.001414668, 0.001413844, 
    0.001410278, 0.001409294, 0.001406578, 0.00140433, 0.001406384, 
    0.001408542, 0.00141467, 0.001420197, 0.001426225, 0.001427701, 
    0.001434752, 0.001429013, 0.001438487, 0.001430433, 0.001444378, 
    0.001419334, 0.001430195, 0.001410525, 0.001412642, 0.001416473, 
    0.001425264, 0.001420516, 0.001426069, 0.001413811, 0.001407459, 
    0.001405815, 0.00140275, 0.001405885, 0.00140563, 0.00140863, 
    0.001407666, 0.001414874, 0.001411001, 0.001422006, 0.001426024, 
    0.001437382, 0.001444351, 0.001451449, 0.001454585, 0.001455539, 
    0.001455938,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3 =
  1.348949e-06, 1.360497e-06, 1.358248e-06, 1.367592e-06, 1.362404e-06, 
    1.368528e-06, 1.351285e-06, 1.360956e-06, 1.354778e-06, 1.349985e-06, 
    1.385818e-06, 1.368008e-06, 1.404436e-06, 1.392987e-06, 1.421834e-06, 
    1.402651e-06, 1.425718e-06, 1.421277e-06, 1.43466e-06, 1.430819e-06, 
    1.448008e-06, 1.436434e-06, 1.456957e-06, 1.445239e-06, 1.447069e-06, 
    1.436052e-06, 1.371582e-06, 1.383595e-06, 1.370872e-06, 1.372582e-06, 
    1.371814e-06, 1.362511e-06, 1.357835e-06, 1.348066e-06, 1.349837e-06, 
    1.357012e-06, 1.37335e-06, 1.367792e-06, 1.381818e-06, 1.3815e-06, 
    1.3972e-06, 1.39011e-06, 1.416631e-06, 1.409067e-06, 1.430979e-06, 
    1.425452e-06, 1.430719e-06, 1.429121e-06, 1.43074e-06, 1.422638e-06, 
    1.426106e-06, 1.418988e-06, 1.391438e-06, 1.399507e-06, 1.375511e-06, 
    1.361184e-06, 1.351708e-06, 1.345005e-06, 1.345951e-06, 1.347757e-06, 
    1.357054e-06, 1.365824e-06, 1.372527e-06, 1.37702e-06, 1.381454e-06, 
    1.394924e-06, 1.402077e-06, 1.418163e-06, 1.415252e-06, 1.420184e-06, 
    1.424903e-06, 1.432844e-06, 1.431535e-06, 1.43504e-06, 1.420052e-06, 
    1.430004e-06, 1.413594e-06, 1.418073e-06, 1.382666e-06, 1.36929e-06, 
    1.363628e-06, 1.358679e-06, 1.346679e-06, 1.35496e-06, 1.351693e-06, 
    1.359472e-06, 1.364427e-06, 1.361975e-06, 1.377143e-06, 1.371236e-06, 
    1.402501e-06, 1.38899e-06, 1.424352e-06, 1.415849e-06, 1.426394e-06, 
    1.421008e-06, 1.430242e-06, 1.42193e-06, 1.436344e-06, 1.439494e-06, 
    1.437341e-06, 1.445616e-06, 1.421469e-06, 1.430718e-06, 1.361907e-06, 
    1.362307e-06, 1.36417e-06, 1.35599e-06, 1.35549e-06, 1.348017e-06, 
    1.354665e-06, 1.357502e-06, 1.364714e-06, 1.36899e-06, 1.37306e-06, 
    1.382032e-06, 1.392088e-06, 1.40621e-06, 1.416399e-06, 1.42325e-06, 
    1.419047e-06, 1.422757e-06, 1.41861e-06, 1.416667e-06, 1.438313e-06, 
    1.426138e-06, 1.444424e-06, 1.443409e-06, 1.435122e-06, 1.443523e-06, 
    1.362587e-06, 1.360287e-06, 1.352318e-06, 1.358552e-06, 1.347204e-06, 
    1.353551e-06, 1.357207e-06, 1.37136e-06, 1.374478e-06, 1.377374e-06, 
    1.383102e-06, 1.390471e-06, 1.403447e-06, 1.414786e-06, 1.425177e-06, 
    1.424414e-06, 1.424682e-06, 1.427009e-06, 1.42125e-06, 1.427955e-06, 
    1.429082e-06, 1.426136e-06, 1.443273e-06, 1.438366e-06, 1.443387e-06, 
    1.440191e-06, 1.361034e-06, 1.364906e-06, 1.362813e-06, 1.36675e-06, 
    1.363976e-06, 1.376334e-06, 1.38005e-06, 1.397504e-06, 1.390326e-06, 
    1.401758e-06, 1.391485e-06, 1.393302e-06, 1.402133e-06, 1.392038e-06, 
    1.41416e-06, 1.399144e-06, 1.427099e-06, 1.412036e-06, 1.428045e-06, 
    1.425131e-06, 1.429957e-06, 1.434288e-06, 1.439744e-06, 1.449841e-06, 
    1.447499e-06, 1.455963e-06, 1.370688e-06, 1.375729e-06, 1.375284e-06, 
    1.380569e-06, 1.384484e-06, 1.392988e-06, 1.406683e-06, 1.401525e-06, 
    1.411001e-06, 1.412908e-06, 1.398513e-06, 1.407343e-06, 1.379107e-06, 
    1.38365e-06, 1.380943e-06, 1.371084e-06, 1.402712e-06, 1.386435e-06, 
    1.416566e-06, 1.407692e-06, 1.433669e-06, 1.420721e-06, 1.446211e-06, 
    1.45718e-06, 1.467538e-06, 1.479694e-06, 1.378484e-06, 1.375054e-06, 
    1.381197e-06, 1.389722e-06, 1.397653e-06, 1.408234e-06, 1.409319e-06, 
    1.411306e-06, 1.41646e-06, 1.420802e-06, 1.411935e-06, 1.421891e-06, 
    1.384706e-06, 1.404129e-06, 1.373757e-06, 1.382868e-06, 1.389217e-06, 
    1.386429e-06, 1.400934e-06, 1.404364e-06, 1.418346e-06, 1.411108e-06, 
    1.454469e-06, 1.435203e-06, 1.488981e-06, 1.473852e-06, 1.373856e-06, 
    1.378471e-06, 1.394595e-06, 1.386911e-06, 1.408941e-06, 1.414391e-06, 
    1.418829e-06, 1.424513e-06, 1.425126e-06, 1.4285e-06, 1.422973e-06, 
    1.428281e-06, 1.408255e-06, 1.417187e-06, 1.392745e-06, 1.398674e-06, 
    1.395945e-06, 1.392954e-06, 1.402194e-06, 1.412073e-06, 1.412283e-06, 
    1.415459e-06, 1.42443e-06, 1.409028e-06, 1.456967e-06, 1.427267e-06, 
    1.383513e-06, 1.392442e-06, 1.393718e-06, 1.390254e-06, 1.413844e-06, 
    1.405273e-06, 1.428418e-06, 1.422143e-06, 1.432431e-06, 1.427314e-06, 
    1.426562e-06, 1.420005e-06, 1.415931e-06, 1.405665e-06, 1.397339e-06, 
    1.390755e-06, 1.392284e-06, 1.399522e-06, 1.412678e-06, 1.425181e-06, 
    1.422437e-06, 1.431646e-06, 1.407335e-06, 1.417504e-06, 1.413569e-06, 
    1.423839e-06, 1.401387e-06, 1.420501e-06, 1.396523e-06, 1.398617e-06, 
    1.405103e-06, 1.418198e-06, 1.421101e-06, 1.424207e-06, 1.42229e-06, 
    1.413014e-06, 1.411496e-06, 1.404944e-06, 1.403138e-06, 1.398159e-06, 
    1.394044e-06, 1.397804e-06, 1.401758e-06, 1.413016e-06, 1.423201e-06, 
    1.434348e-06, 1.437082e-06, 1.450177e-06, 1.439514e-06, 1.457133e-06, 
    1.442149e-06, 1.468135e-06, 1.42161e-06, 1.44171e-06, 1.405398e-06, 
    1.409287e-06, 1.416336e-06, 1.432569e-06, 1.423792e-06, 1.434059e-06, 
    1.411437e-06, 1.399773e-06, 1.396761e-06, 1.391154e-06, 1.396889e-06, 
    1.396422e-06, 1.401921e-06, 1.400152e-06, 1.41339e-06, 1.406271e-06, 
    1.426541e-06, 1.433975e-06, 1.455073e-06, 1.468085e-06, 1.481388e-06, 
    1.487281e-06, 1.489077e-06, 1.489828e-06 ;

 SMIN_NO3_LEACHED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_RUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_vr =
  8.30805e-06, 8.344628e-06, 8.337495e-06, 8.367022e-06, 8.350627e-06, 
    8.369953e-06, 8.315418e-06, 8.34603e-06, 8.326471e-06, 8.311266e-06, 
    8.424324e-06, 8.368273e-06, 8.482571e-06, 8.446762e-06, 8.536713e-06, 
    8.476982e-06, 8.548755e-06, 8.534957e-06, 8.576433e-06, 8.564532e-06, 
    8.617637e-06, 8.581898e-06, 8.645161e-06, 8.609079e-06, 8.614716e-06, 
    8.580681e-06, 8.379596e-06, 8.417405e-06, 8.377343e-06, 8.382734e-06, 
    8.380302e-06, 8.350934e-06, 8.336152e-06, 8.305175e-06, 8.310782e-06, 
    8.333524e-06, 8.385097e-06, 8.36756e-06, 8.411709e-06, 8.410713e-06, 
    8.459914e-06, 8.437718e-06, 8.520507e-06, 8.496943e-06, 8.565019e-06, 
    8.547878e-06, 8.5642e-06, 8.559235e-06, 8.56424e-06, 8.539123e-06, 
    8.549866e-06, 8.527767e-06, 8.441973e-06, 8.467214e-06, 8.39194e-06, 
    8.346746e-06, 8.316728e-06, 8.295457e-06, 8.298446e-06, 8.304182e-06, 
    8.333641e-06, 8.361346e-06, 8.38248e-06, 8.396614e-06, 8.410546e-06, 
    8.452802e-06, 8.47515e-06, 8.525257e-06, 8.516196e-06, 8.531521e-06, 
    8.546164e-06, 8.570762e-06, 8.566706e-06, 8.577541e-06, 8.531067e-06, 
    8.561947e-06, 8.510968e-06, 8.524903e-06, 8.414453e-06, 8.372323e-06, 
    8.354459e-06, 8.338793e-06, 8.300753e-06, 8.327016e-06, 8.316651e-06, 
    8.341268e-06, 8.356926e-06, 8.349165e-06, 8.396993e-06, 8.378379e-06, 
    8.476462e-06, 8.434185e-06, 8.544466e-06, 8.518035e-06, 8.550775e-06, 
    8.534061e-06, 8.562692e-06, 8.536908e-06, 8.58156e-06, 8.591297e-06, 
    8.584627e-06, 8.610178e-06, 8.53543e-06, 8.564121e-06, 8.348998e-06, 
    8.350263e-06, 8.356137e-06, 8.330265e-06, 8.328679e-06, 8.304973e-06, 
    8.32604e-06, 8.335024e-06, 8.35781e-06, 8.371293e-06, 8.384113e-06, 
    8.41234e-06, 8.443877e-06, 8.488008e-06, 8.519739e-06, 8.541012e-06, 
    8.527953e-06, 8.539467e-06, 8.526579e-06, 8.520527e-06, 8.587627e-06, 
    8.549937e-06, 8.606478e-06, 8.603347e-06, 8.577736e-06, 8.603676e-06, 
    8.351134e-06, 8.34385e-06, 8.318622e-06, 8.338348e-06, 8.302377e-06, 
    8.322509e-06, 8.334078e-06, 8.378764e-06, 8.388572e-06, 8.397691e-06, 
    8.415685e-06, 8.438791e-06, 8.479377e-06, 8.514705e-06, 8.546981e-06, 
    8.544602e-06, 8.545432e-06, 8.552636e-06, 8.534761e-06, 8.555555e-06, 
    8.55904e-06, 8.549907e-06, 8.602904e-06, 8.587754e-06, 8.603248e-06, 
    8.593367e-06, 8.346203e-06, 8.358425e-06, 8.351803e-06, 8.36424e-06, 
    8.355464e-06, 8.394431e-06, 8.40611e-06, 8.460825e-06, 8.438337e-06, 
    8.474109e-06, 8.441951e-06, 8.447648e-06, 8.475263e-06, 8.443663e-06, 
    8.512737e-06, 8.465893e-06, 8.552908e-06, 8.506103e-06, 8.555826e-06, 
    8.546775e-06, 8.561727e-06, 8.575138e-06, 8.591987e-06, 8.623139e-06, 
    8.615904e-06, 8.641962e-06, 8.376658e-06, 8.39253e-06, 8.391122e-06, 
    8.407733e-06, 8.420022e-06, 8.446686e-06, 8.489478e-06, 8.473363e-06, 
    8.502911e-06, 8.508852e-06, 8.463924e-06, 8.491501e-06, 8.403074e-06, 
    8.417342e-06, 8.408831e-06, 8.37779e-06, 8.477014e-06, 8.426054e-06, 
    8.520166e-06, 8.49252e-06, 8.573203e-06, 8.533062e-06, 8.611928e-06, 
    8.645708e-06, 8.677477e-06, 8.714662e-06, 8.401185e-06, 8.390378e-06, 
    8.409692e-06, 8.436456e-06, 8.461265e-06, 8.494305e-06, 8.497672e-06, 
    8.503854e-06, 8.519883e-06, 8.53338e-06, 8.505798e-06, 8.536739e-06, 
    8.420658e-06, 8.481434e-06, 8.386196e-06, 8.414861e-06, 8.43476e-06, 
    8.426017e-06, 8.471415e-06, 8.482113e-06, 8.525657e-06, 8.503135e-06, 
    8.63735e-06, 8.577918e-06, 8.742964e-06, 8.69679e-06, 8.386599e-06, 
    8.401111e-06, 8.451695e-06, 8.427615e-06, 8.496483e-06, 8.51346e-06, 
    8.52724e-06, 8.544897e-06, 8.546781e-06, 8.557246e-06, 8.540084e-06, 
    8.556551e-06, 8.494286e-06, 8.522094e-06, 8.445812e-06, 8.464354e-06, 
    8.455811e-06, 8.446438e-06, 8.475324e-06, 8.506142e-06, 8.50678e-06, 
    8.516654e-06, 8.544542e-06, 8.496611e-06, 8.645015e-06, 8.553312e-06, 
    8.416945e-06, 8.444946e-06, 8.448925e-06, 8.438074e-06, 8.511735e-06, 
    8.485028e-06, 8.55699e-06, 8.537512e-06, 8.569396e-06, 8.553547e-06, 
    8.551197e-06, 8.530847e-06, 8.518166e-06, 8.486189e-06, 8.460165e-06, 
    8.43955e-06, 8.444325e-06, 8.466976e-06, 8.508001e-06, 8.546856e-06, 
    8.538334e-06, 8.566868e-06, 8.491317e-06, 8.522985e-06, 8.510729e-06, 
    8.542645e-06, 8.472904e-06, 8.532465e-06, 8.457687e-06, 8.464222e-06, 
    8.484473e-06, 8.525265e-06, 8.53426e-06, 8.543907e-06, 8.537935e-06, 
    8.509102e-06, 8.504365e-06, 8.483925e-06, 8.478281e-06, 8.462723e-06, 
    8.449831e-06, 8.461598e-06, 8.473939e-06, 8.509046e-06, 8.540698e-06, 
    8.575229e-06, 8.583678e-06, 8.624089e-06, 8.591191e-06, 8.645487e-06, 
    8.599327e-06, 8.679228e-06, 8.535879e-06, 8.598119e-06, 8.485394e-06, 
    8.497509e-06, 8.519459e-06, 8.569818e-06, 8.542595e-06, 8.574417e-06, 
    8.504174e-06, 8.467776e-06, 8.458343e-06, 8.440794e-06, 8.458729e-06, 
    8.45727e-06, 8.474445e-06, 8.468909e-06, 8.510187e-06, 8.488006e-06, 
    8.551033e-06, 8.574065e-06, 8.639139e-06, 8.679074e-06, 8.719749e-06, 
    8.737709e-06, 8.743176e-06, 8.745455e-06,
  4.946847e-06, 4.984e-06, 4.976769e-06, 5.006795e-06, 4.99013e-06, 
    5.009803e-06, 4.95437e-06, 4.985479e-06, 4.965611e-06, 4.950185e-06, 
    5.065255e-06, 5.008136e-06, 5.124812e-06, 5.088208e-06, 5.180328e-06, 
    5.119112e-06, 5.192701e-06, 5.178554e-06, 5.221164e-06, 5.208944e-06, 
    5.263584e-06, 5.226806e-06, 5.291979e-06, 5.254791e-06, 5.260604e-06, 
    5.225595e-06, 5.019608e-06, 5.058133e-06, 5.01733e-06, 5.022816e-06, 
    5.020353e-06, 4.990475e-06, 4.975445e-06, 4.944008e-06, 4.949709e-06, 
    4.9728e-06, 5.025283e-06, 5.007443e-06, 5.052441e-06, 5.051423e-06, 
    5.101685e-06, 5.079001e-06, 5.163741e-06, 5.139605e-06, 5.209454e-06, 
    5.191857e-06, 5.208627e-06, 5.20354e-06, 5.208693e-06, 5.182895e-06, 
    5.193943e-06, 5.17126e-06, 5.083248e-06, 5.109061e-06, 5.032215e-06, 
    4.986213e-06, 4.955733e-06, 4.934148e-06, 4.937197e-06, 4.943014e-06, 
    4.972935e-06, 5.001124e-06, 5.022645e-06, 5.03706e-06, 5.051277e-06, 
    5.094408e-06, 5.117279e-06, 5.168628e-06, 5.159344e-06, 5.175072e-06, 
    5.190107e-06, 5.215391e-06, 5.211225e-06, 5.222375e-06, 5.174654e-06, 
    5.206354e-06, 5.15406e-06, 5.168345e-06, 5.055158e-06, 5.012253e-06, 
    4.994068e-06, 4.978159e-06, 4.939543e-06, 4.9662e-06, 4.955686e-06, 
    4.98071e-06, 4.996636e-06, 4.988756e-06, 5.037454e-06, 5.018502e-06, 
    5.118636e-06, 5.075419e-06, 5.188353e-06, 5.161249e-06, 5.194857e-06, 
    5.177697e-06, 5.207112e-06, 5.180636e-06, 5.226526e-06, 5.236539e-06, 
    5.229696e-06, 5.255994e-06, 5.17917e-06, 5.208628e-06, 4.988536e-06, 
    4.989821e-06, 4.995808e-06, 4.969514e-06, 4.967906e-06, 4.943853e-06, 
    4.965252e-06, 4.974376e-06, 4.997559e-06, 5.011292e-06, 5.024359e-06, 
    5.053131e-06, 5.085335e-06, 5.130484e-06, 5.163005e-06, 5.184845e-06, 
    5.171448e-06, 5.183275e-06, 5.170054e-06, 5.163862e-06, 5.232787e-06, 
    5.194047e-06, 5.252208e-06, 5.248984e-06, 5.222641e-06, 5.249347e-06, 
    4.990723e-06, 4.983331e-06, 4.9577e-06, 4.977754e-06, 4.941236e-06, 
    4.961667e-06, 4.973429e-06, 5.018901e-06, 5.028908e-06, 5.038198e-06, 
    5.05656e-06, 5.080162e-06, 5.121659e-06, 5.15786e-06, 5.190982e-06, 
    5.188553e-06, 5.189408e-06, 5.196818e-06, 5.178471e-06, 5.199832e-06, 
    5.203422e-06, 5.194041e-06, 5.248552e-06, 5.232958e-06, 5.248915e-06, 
    5.23876e-06, 4.985733e-06, 4.998175e-06, 4.991451e-06, 5.0041e-06, 
    4.995188e-06, 5.03486e-06, 5.046777e-06, 5.102664e-06, 5.079698e-06, 
    5.116261e-06, 5.083406e-06, 5.089224e-06, 5.117462e-06, 5.085179e-06, 
    5.155865e-06, 5.10791e-06, 5.197106e-06, 5.14909e-06, 5.200121e-06, 
    5.190839e-06, 5.206208e-06, 5.219988e-06, 5.237339e-06, 5.26941e-06, 
    5.261977e-06, 5.288834e-06, 5.016744e-06, 5.032922e-06, 5.031494e-06, 
    5.048441e-06, 5.060987e-06, 5.088215e-06, 5.131997e-06, 5.115517e-06, 
    5.145783e-06, 5.151867e-06, 5.10589e-06, 5.134105e-06, 5.043757e-06, 
    5.058319e-06, 5.049646e-06, 5.018021e-06, 5.119316e-06, 5.067243e-06, 
    5.163543e-06, 5.135224e-06, 5.218023e-06, 5.176791e-06, 5.257888e-06, 
    5.292695e-06, 5.325513e-06, 5.363966e-06, 5.041757e-06, 5.030755e-06, 
    5.050457e-06, 5.077764e-06, 5.103141e-06, 5.136951e-06, 5.140413e-06, 
    5.146758e-06, 5.163202e-06, 5.177044e-06, 5.148767e-06, 5.180515e-06, 
    5.061703e-06, 5.123844e-06, 5.0266e-06, 5.055817e-06, 5.076152e-06, 
    5.067226e-06, 5.113634e-06, 5.124594e-06, 5.16922e-06, 5.146132e-06, 
    5.2841e-06, 5.222904e-06, 5.393298e-06, 5.345496e-06, 5.026914e-06, 
    5.041717e-06, 5.09336e-06, 5.068765e-06, 5.139209e-06, 5.156602e-06, 
    5.170754e-06, 5.188869e-06, 5.190824e-06, 5.201568e-06, 5.183966e-06, 
    5.200872e-06, 5.137023e-06, 5.165521e-06, 5.087445e-06, 5.106411e-06, 
    5.097682e-06, 5.088115e-06, 5.117663e-06, 5.149212e-06, 5.149883e-06, 
    5.160015e-06, 5.188612e-06, 5.139495e-06, 5.292024e-06, 5.197651e-06, 
    5.057877e-06, 5.086471e-06, 5.090555e-06, 5.079469e-06, 5.154858e-06, 
    5.127497e-06, 5.201306e-06, 5.181321e-06, 5.214079e-06, 5.197792e-06, 
    5.195398e-06, 5.174508e-06, 5.161519e-06, 5.128751e-06, 5.102143e-06, 
    5.081076e-06, 5.085972e-06, 5.109123e-06, 5.151143e-06, 5.191003e-06, 
    5.182263e-06, 5.211587e-06, 5.13409e-06, 5.166539e-06, 5.15399e-06, 
    5.186732e-06, 5.11508e-06, 5.176087e-06, 5.099529e-06, 5.106224e-06, 
    5.126954e-06, 5.168745e-06, 5.178e-06, 5.187897e-06, 5.181789e-06, 
    5.152211e-06, 5.147369e-06, 5.126449e-06, 5.120681e-06, 5.104765e-06, 
    5.091605e-06, 5.10363e-06, 5.11627e-06, 5.152222e-06, 5.184698e-06, 
    5.220185e-06, 5.228881e-06, 5.270484e-06, 5.236614e-06, 5.292552e-06, 
    5.24499e-06, 5.327409e-06, 5.179623e-06, 5.243585e-06, 5.127897e-06, 
    5.140316e-06, 5.16281e-06, 5.214521e-06, 5.186577e-06, 5.219261e-06, 
    5.147179e-06, 5.109924e-06, 5.100296e-06, 5.082357e-06, 5.100706e-06, 
    5.099213e-06, 5.116791e-06, 5.11114e-06, 5.153417e-06, 5.130692e-06, 
    5.195339e-06, 5.219001e-06, 5.286019e-06, 5.32725e-06, 5.369324e-06, 
    5.387936e-06, 5.393605e-06, 5.395976e-06,
  4.461329e-06, 4.500614e-06, 4.492965e-06, 4.524734e-06, 4.507098e-06, 
    4.527918e-06, 4.469281e-06, 4.502177e-06, 4.481165e-06, 4.464858e-06, 
    4.586655e-06, 4.526153e-06, 4.649839e-06, 4.610998e-06, 4.708818e-06, 
    4.643787e-06, 4.721975e-06, 4.706934e-06, 4.752256e-06, 4.739254e-06, 
    4.797421e-06, 4.758262e-06, 4.827682e-06, 4.788056e-06, 4.794248e-06, 
    4.756972e-06, 4.538299e-06, 4.579105e-06, 4.535887e-06, 4.541695e-06, 
    4.539088e-06, 4.507463e-06, 4.491563e-06, 4.45833e-06, 4.464356e-06, 
    4.488767e-06, 4.544308e-06, 4.525421e-06, 4.573079e-06, 4.572e-06, 
    4.625295e-06, 4.601234e-06, 4.691189e-06, 4.665549e-06, 4.739796e-06, 
    4.721079e-06, 4.738917e-06, 4.733505e-06, 4.738987e-06, 4.711549e-06, 
    4.723297e-06, 4.699181e-06, 4.605737e-06, 4.633121e-06, 4.551649e-06, 
    4.502952e-06, 4.470722e-06, 4.447911e-06, 4.451133e-06, 4.457278e-06, 
    4.48891e-06, 4.518733e-06, 4.541515e-06, 4.556782e-06, 4.571845e-06, 
    4.617571e-06, 4.641842e-06, 4.696382e-06, 4.686518e-06, 4.703232e-06, 
    4.719218e-06, 4.746112e-06, 4.741681e-06, 4.753545e-06, 4.702789e-06, 
    4.736498e-06, 4.680903e-06, 4.696083e-06, 4.575953e-06, 4.530512e-06, 
    4.511263e-06, 4.494435e-06, 4.453611e-06, 4.481788e-06, 4.470671e-06, 
    4.497134e-06, 4.513983e-06, 4.505646e-06, 4.5572e-06, 4.537128e-06, 
    4.643282e-06, 4.597434e-06, 4.717353e-06, 4.688542e-06, 4.724269e-06, 
    4.706024e-06, 4.737304e-06, 4.709148e-06, 4.757963e-06, 4.76862e-06, 
    4.761337e-06, 4.789338e-06, 4.70759e-06, 4.738918e-06, 4.505413e-06, 
    4.506772e-06, 4.513106e-06, 4.485291e-06, 4.483592e-06, 4.458166e-06, 
    4.480786e-06, 4.490434e-06, 4.51496e-06, 4.529495e-06, 4.54333e-06, 
    4.573809e-06, 4.607949e-06, 4.655862e-06, 4.690407e-06, 4.713622e-06, 
    4.699381e-06, 4.711953e-06, 4.6979e-06, 4.691319e-06, 4.764627e-06, 
    4.723407e-06, 4.785306e-06, 4.781873e-06, 4.753828e-06, 4.78226e-06, 
    4.507727e-06, 4.499906e-06, 4.472801e-06, 4.494007e-06, 4.4554e-06, 
    4.476995e-06, 4.489432e-06, 4.53755e-06, 4.548148e-06, 4.557987e-06, 
    4.577444e-06, 4.602464e-06, 4.646493e-06, 4.68494e-06, 4.720149e-06, 
    4.717565e-06, 4.718475e-06, 4.726355e-06, 4.706847e-06, 4.729561e-06, 
    4.733378e-06, 4.723401e-06, 4.781413e-06, 4.76481e-06, 4.781799e-06, 
    4.770986e-06, 4.502448e-06, 4.515613e-06, 4.508497e-06, 4.521882e-06, 
    4.512451e-06, 4.554451e-06, 4.567074e-06, 4.626332e-06, 4.601972e-06, 
    4.640763e-06, 4.605905e-06, 4.612074e-06, 4.642035e-06, 4.607786e-06, 
    4.682819e-06, 4.631898e-06, 4.726662e-06, 4.67562e-06, 4.729868e-06, 
    4.719996e-06, 4.736343e-06, 4.751005e-06, 4.769473e-06, 4.80363e-06, 
    4.795711e-06, 4.824332e-06, 4.535267e-06, 4.552398e-06, 4.550887e-06, 
    4.568839e-06, 4.582135e-06, 4.611006e-06, 4.657469e-06, 4.639974e-06, 
    4.67211e-06, 4.678574e-06, 4.629757e-06, 4.659707e-06, 4.563877e-06, 
    4.579306e-06, 4.570115e-06, 4.536619e-06, 4.644005e-06, 4.588766e-06, 
    4.690979e-06, 4.660896e-06, 4.748913e-06, 4.705058e-06, 4.791355e-06, 
    4.828445e-06, 4.863449e-06, 4.904494e-06, 4.561757e-06, 4.550104e-06, 
    4.570976e-06, 4.599921e-06, 4.626839e-06, 4.662729e-06, 4.666407e-06, 
    4.673146e-06, 4.690618e-06, 4.705329e-06, 4.675279e-06, 4.70902e-06, 
    4.58289e-06, 4.648812e-06, 4.545703e-06, 4.576654e-06, 4.598211e-06, 
    4.588748e-06, 4.637976e-06, 4.64961e-06, 4.697011e-06, 4.672482e-06, 
    4.819282e-06, 4.754106e-06, 4.935832e-06, 4.884773e-06, 4.546036e-06, 
    4.561716e-06, 4.616463e-06, 4.59038e-06, 4.665128e-06, 4.683604e-06, 
    4.698644e-06, 4.717901e-06, 4.719981e-06, 4.731407e-06, 4.712689e-06, 
    4.730667e-06, 4.662806e-06, 4.693082e-06, 4.610189e-06, 4.63031e-06, 
    4.621048e-06, 4.6109e-06, 4.642251e-06, 4.675752e-06, 4.676466e-06, 
    4.68723e-06, 4.717622e-06, 4.665432e-06, 4.827726e-06, 4.727235e-06, 
    4.578839e-06, 4.609154e-06, 4.613487e-06, 4.60173e-06, 4.68175e-06, 
    4.652691e-06, 4.731128e-06, 4.709876e-06, 4.744717e-06, 4.727391e-06, 
    4.724845e-06, 4.702634e-06, 4.688829e-06, 4.654023e-06, 4.625781e-06, 
    4.603435e-06, 4.608627e-06, 4.633187e-06, 4.677804e-06, 4.72017e-06, 
    4.710877e-06, 4.742065e-06, 4.659692e-06, 4.694162e-06, 4.680828e-06, 
    4.715629e-06, 4.63951e-06, 4.704306e-06, 4.623007e-06, 4.630112e-06, 
    4.652115e-06, 4.696506e-06, 4.706346e-06, 4.716867e-06, 4.710374e-06, 
    4.678938e-06, 4.673795e-06, 4.651579e-06, 4.645454e-06, 4.628565e-06, 
    4.614601e-06, 4.627359e-06, 4.640773e-06, 4.67895e-06, 4.713466e-06, 
    4.751214e-06, 4.760469e-06, 4.804771e-06, 4.768699e-06, 4.828288e-06, 
    4.777613e-06, 4.865467e-06, 4.708068e-06, 4.77612e-06, 4.653116e-06, 
    4.666304e-06, 4.690199e-06, 4.745186e-06, 4.715465e-06, 4.750229e-06, 
    4.673593e-06, 4.634036e-06, 4.623821e-06, 4.604792e-06, 4.624257e-06, 
    4.622672e-06, 4.641327e-06, 4.635328e-06, 4.68022e-06, 4.656084e-06, 
    4.724781e-06, 4.749953e-06, 4.82133e-06, 4.865301e-06, 4.910219e-06, 
    4.930103e-06, 4.936162e-06, 4.938695e-06,
  4.331477e-06, 4.372477e-06, 4.364491e-06, 4.397667e-06, 4.379247e-06, 
    4.400993e-06, 4.339774e-06, 4.37411e-06, 4.352175e-06, 4.335159e-06, 
    4.46239e-06, 4.399149e-06, 4.528519e-06, 4.487857e-06, 4.590327e-06, 
    4.522182e-06, 4.604125e-06, 4.58835e-06, 4.635895e-06, 4.62225e-06, 
    4.683322e-06, 4.642198e-06, 4.715122e-06, 4.673483e-06, 4.679987e-06, 
    4.640845e-06, 4.411838e-06, 4.454495e-06, 4.409318e-06, 4.415387e-06, 
    4.412662e-06, 4.379629e-06, 4.363028e-06, 4.328349e-06, 4.334635e-06, 
    4.360109e-06, 4.418117e-06, 4.398383e-06, 4.448191e-06, 4.447063e-06, 
    4.502821e-06, 4.47764e-06, 4.571844e-06, 4.544975e-06, 4.62282e-06, 
    4.603184e-06, 4.621897e-06, 4.616219e-06, 4.621971e-06, 4.593189e-06, 
    4.605511e-06, 4.580222e-06, 4.482352e-06, 4.511013e-06, 4.425789e-06, 
    4.374919e-06, 4.341277e-06, 4.317481e-06, 4.320842e-06, 4.327252e-06, 
    4.360259e-06, 4.391397e-06, 4.415198e-06, 4.431154e-06, 4.446901e-06, 
    4.494736e-06, 4.520145e-06, 4.577288e-06, 4.566948e-06, 4.584469e-06, 
    4.601233e-06, 4.629447e-06, 4.624797e-06, 4.637248e-06, 4.584004e-06, 
    4.619359e-06, 4.561063e-06, 4.576973e-06, 4.451198e-06, 4.403702e-06, 
    4.383597e-06, 4.366026e-06, 4.323426e-06, 4.352825e-06, 4.341225e-06, 
    4.368843e-06, 4.386437e-06, 4.377731e-06, 4.431591e-06, 4.410615e-06, 
    4.521653e-06, 4.473665e-06, 4.599276e-06, 4.569069e-06, 4.60653e-06, 
    4.587396e-06, 4.620205e-06, 4.590672e-06, 4.641885e-06, 4.653074e-06, 
    4.645427e-06, 4.67483e-06, 4.589038e-06, 4.621898e-06, 4.377488e-06, 
    4.378907e-06, 4.385522e-06, 4.356482e-06, 4.354707e-06, 4.328178e-06, 
    4.351779e-06, 4.361849e-06, 4.387457e-06, 4.40264e-06, 4.417095e-06, 
    4.448955e-06, 4.484667e-06, 4.534827e-06, 4.571024e-06, 4.595364e-06, 
    4.580431e-06, 4.593614e-06, 4.578879e-06, 4.571979e-06, 4.648881e-06, 
    4.605626e-06, 4.670595e-06, 4.666988e-06, 4.637545e-06, 4.667395e-06, 
    4.379904e-06, 4.371738e-06, 4.343447e-06, 4.36558e-06, 4.325293e-06, 
    4.347823e-06, 4.360804e-06, 4.411055e-06, 4.42213e-06, 4.432414e-06, 
    4.452756e-06, 4.478928e-06, 4.525015e-06, 4.565294e-06, 4.602209e-06, 
    4.599499e-06, 4.600453e-06, 4.608718e-06, 4.588259e-06, 4.612081e-06, 
    4.616086e-06, 4.60562e-06, 4.666505e-06, 4.649073e-06, 4.666912e-06, 
    4.655557e-06, 4.374391e-06, 4.388139e-06, 4.380708e-06, 4.394687e-06, 
    4.384837e-06, 4.428718e-06, 4.441914e-06, 4.503906e-06, 4.478412e-06, 
    4.519015e-06, 4.482528e-06, 4.488984e-06, 4.520347e-06, 4.484496e-06, 
    4.563071e-06, 4.509733e-06, 4.60904e-06, 4.555528e-06, 4.612403e-06, 
    4.602049e-06, 4.619197e-06, 4.634582e-06, 4.653969e-06, 4.689844e-06, 
    4.681525e-06, 4.711599e-06, 4.40867e-06, 4.426572e-06, 4.424992e-06, 
    4.443759e-06, 4.457663e-06, 4.487865e-06, 4.53651e-06, 4.518188e-06, 
    4.551849e-06, 4.558622e-06, 4.507491e-06, 4.538855e-06, 4.438571e-06, 
    4.454704e-06, 4.445093e-06, 4.410082e-06, 4.52241e-06, 4.464598e-06, 
    4.571624e-06, 4.540101e-06, 4.632387e-06, 4.586384e-06, 4.676948e-06, 
    4.715924e-06, 4.752733e-06, 4.795932e-06, 4.436355e-06, 4.424174e-06, 
    4.445993e-06, 4.476267e-06, 4.504437e-06, 4.542021e-06, 4.545873e-06, 
    4.552934e-06, 4.571245e-06, 4.586668e-06, 4.55517e-06, 4.590538e-06, 
    4.458453e-06, 4.527444e-06, 4.419575e-06, 4.451931e-06, 4.474479e-06, 
    4.464579e-06, 4.516095e-06, 4.528279e-06, 4.577947e-06, 4.552238e-06, 
    4.706292e-06, 4.637838e-06, 4.828938e-06, 4.775171e-06, 4.419923e-06, 
    4.436311e-06, 4.493576e-06, 4.466286e-06, 4.544534e-06, 4.563894e-06, 
    4.579658e-06, 4.599851e-06, 4.602032e-06, 4.614019e-06, 4.594385e-06, 
    4.613241e-06, 4.542101e-06, 4.573827e-06, 4.48701e-06, 4.50807e-06, 
    4.498375e-06, 4.487754e-06, 4.520573e-06, 4.555665e-06, 4.556413e-06, 
    4.567694e-06, 4.59956e-06, 4.544852e-06, 4.715168e-06, 4.609644e-06, 
    4.454215e-06, 4.485928e-06, 4.490462e-06, 4.47816e-06, 4.561951e-06, 
    4.531506e-06, 4.613726e-06, 4.591435e-06, 4.627983e-06, 4.609805e-06, 
    4.607134e-06, 4.583841e-06, 4.569369e-06, 4.532901e-06, 4.503329e-06, 
    4.479943e-06, 4.485375e-06, 4.511082e-06, 4.557815e-06, 4.602231e-06, 
    4.592485e-06, 4.625201e-06, 4.538839e-06, 4.574961e-06, 4.560985e-06, 
    4.597468e-06, 4.517702e-06, 4.585597e-06, 4.500426e-06, 4.507863e-06, 
    4.530903e-06, 4.577418e-06, 4.587734e-06, 4.598767e-06, 4.591957e-06, 
    4.559004e-06, 4.553614e-06, 4.530341e-06, 4.523928e-06, 4.506242e-06, 
    4.491628e-06, 4.504981e-06, 4.519025e-06, 4.559016e-06, 4.5952e-06, 
    4.634802e-06, 4.644516e-06, 4.691044e-06, 4.653157e-06, 4.71576e-06, 
    4.662518e-06, 4.754858e-06, 4.58954e-06, 4.660949e-06, 4.531951e-06, 
    4.545766e-06, 4.570807e-06, 4.628476e-06, 4.597296e-06, 4.633769e-06, 
    4.553403e-06, 4.511972e-06, 4.501278e-06, 4.481363e-06, 4.501733e-06, 
    4.500075e-06, 4.519604e-06, 4.513324e-06, 4.560347e-06, 4.535059e-06, 
    4.607068e-06, 4.633479e-06, 4.708444e-06, 4.754681e-06, 4.801959e-06, 
    4.822903e-06, 4.829285e-06, 4.831955e-06,
  4.364439e-06, 4.40508e-06, 4.397161e-06, 4.430066e-06, 4.411794e-06, 
    4.433366e-06, 4.372659e-06, 4.4067e-06, 4.38495e-06, 4.368086e-06, 
    4.494324e-06, 4.431537e-06, 4.56006e-06, 4.519628e-06, 4.621583e-06, 
    4.553758e-06, 4.635328e-06, 4.619614e-06, 4.666991e-06, 4.653389e-06, 
    4.714299e-06, 4.673276e-06, 4.746046e-06, 4.704481e-06, 4.710972e-06, 
    4.671926e-06, 4.444128e-06, 4.486481e-06, 4.441627e-06, 4.44765e-06, 
    4.444946e-06, 4.412173e-06, 4.395712e-06, 4.361338e-06, 4.367566e-06, 
    4.392817e-06, 4.45036e-06, 4.430776e-06, 4.480218e-06, 4.479098e-06, 
    4.534503e-06, 4.509474e-06, 4.603176e-06, 4.576431e-06, 4.653956e-06, 
    4.63439e-06, 4.653037e-06, 4.647378e-06, 4.653111e-06, 4.624434e-06, 
    4.636708e-06, 4.611518e-06, 4.514156e-06, 4.542649e-06, 4.457975e-06, 
    4.407504e-06, 4.37415e-06, 4.350572e-06, 4.3539e-06, 4.360251e-06, 
    4.392965e-06, 4.423845e-06, 4.447462e-06, 4.463301e-06, 4.478937e-06, 
    4.526468e-06, 4.551731e-06, 4.608597e-06, 4.598301e-06, 4.615748e-06, 
    4.632446e-06, 4.660563e-06, 4.655928e-06, 4.66834e-06, 4.615285e-06, 
    4.650508e-06, 4.592443e-06, 4.608284e-06, 4.483208e-06, 4.436054e-06, 
    4.41611e-06, 4.398683e-06, 4.356461e-06, 4.385595e-06, 4.374097e-06, 
    4.401476e-06, 4.418926e-06, 4.41029e-06, 4.463734e-06, 4.442913e-06, 
    4.553231e-06, 4.505524e-06, 4.630497e-06, 4.600413e-06, 4.637724e-06, 
    4.618663e-06, 4.651351e-06, 4.621926e-06, 4.672963e-06, 4.684121e-06, 
    4.676495e-06, 4.705824e-06, 4.620298e-06, 4.653039e-06, 4.410048e-06, 
    4.411456e-06, 4.418017e-06, 4.389221e-06, 4.387462e-06, 4.361168e-06, 
    4.384558e-06, 4.394542e-06, 4.419937e-06, 4.435e-06, 4.449344e-06, 
    4.480977e-06, 4.516458e-06, 4.566336e-06, 4.60236e-06, 4.626599e-06, 
    4.611727e-06, 4.624856e-06, 4.610181e-06, 4.603311e-06, 4.67994e-06, 
    4.636824e-06, 4.701599e-06, 4.698001e-06, 4.668636e-06, 4.698406e-06, 
    4.412445e-06, 4.404346e-06, 4.3763e-06, 4.39824e-06, 4.35831e-06, 
    4.380638e-06, 4.393506e-06, 4.443351e-06, 4.454342e-06, 4.464552e-06, 
    4.484752e-06, 4.510753e-06, 4.556574e-06, 4.596656e-06, 4.633418e-06, 
    4.630719e-06, 4.631669e-06, 4.639904e-06, 4.619522e-06, 4.643255e-06, 
    4.647246e-06, 4.636817e-06, 4.697519e-06, 4.68013e-06, 4.697924e-06, 
    4.686597e-06, 4.406977e-06, 4.420613e-06, 4.413242e-06, 4.427109e-06, 
    4.417338e-06, 4.460883e-06, 4.473985e-06, 4.535583e-06, 4.510242e-06, 
    4.550607e-06, 4.514331e-06, 4.520748e-06, 4.551933e-06, 4.516286e-06, 
    4.594443e-06, 4.541377e-06, 4.640224e-06, 4.586936e-06, 4.643576e-06, 
    4.633259e-06, 4.650346e-06, 4.665682e-06, 4.685014e-06, 4.720809e-06, 
    4.712505e-06, 4.742528e-06, 4.440984e-06, 4.458752e-06, 4.457184e-06, 
    4.475817e-06, 4.489626e-06, 4.519636e-06, 4.568009e-06, 4.549784e-06, 
    4.583273e-06, 4.590013e-06, 4.539146e-06, 4.570342e-06, 4.470665e-06, 
    4.486687e-06, 4.477142e-06, 4.442385e-06, 4.553984e-06, 4.496516e-06, 
    4.602957e-06, 4.571581e-06, 4.663494e-06, 4.617656e-06, 4.707938e-06, 
    4.746848e-06, 4.783622e-06, 4.826822e-06, 4.468464e-06, 4.456371e-06, 
    4.478034e-06, 4.50811e-06, 4.53611e-06, 4.573492e-06, 4.577325e-06, 
    4.584353e-06, 4.602579e-06, 4.617938e-06, 4.586578e-06, 4.621792e-06, 
    4.490413e-06, 4.55899e-06, 4.451807e-06, 4.483933e-06, 4.506333e-06, 
    4.496496e-06, 4.547702e-06, 4.55982e-06, 4.609254e-06, 4.58366e-06, 
    4.73723e-06, 4.668929e-06, 4.859856e-06, 4.806057e-06, 4.452151e-06, 
    4.468421e-06, 4.525313e-06, 4.498192e-06, 4.575993e-06, 4.595261e-06, 
    4.610957e-06, 4.63107e-06, 4.633242e-06, 4.645186e-06, 4.625624e-06, 
    4.644411e-06, 4.573572e-06, 4.605151e-06, 4.518786e-06, 4.539722e-06, 
    4.530083e-06, 4.519525e-06, 4.552156e-06, 4.587072e-06, 4.587815e-06, 
    4.599045e-06, 4.630783e-06, 4.576309e-06, 4.746096e-06, 4.640829e-06, 
    4.486201e-06, 4.517712e-06, 4.522217e-06, 4.50999e-06, 4.593328e-06, 
    4.563031e-06, 4.644894e-06, 4.622686e-06, 4.659104e-06, 4.640987e-06, 
    4.638325e-06, 4.615123e-06, 4.600713e-06, 4.564419e-06, 4.535008e-06, 
    4.511761e-06, 4.517161e-06, 4.542718e-06, 4.589212e-06, 4.633441e-06, 
    4.623732e-06, 4.65633e-06, 4.570326e-06, 4.60628e-06, 4.592366e-06, 
    4.628695e-06, 4.549301e-06, 4.616874e-06, 4.532122e-06, 4.539515e-06, 
    4.562431e-06, 4.608728e-06, 4.618999e-06, 4.62999e-06, 4.623205e-06, 
    4.590394e-06, 4.58503e-06, 4.561872e-06, 4.555493e-06, 4.537905e-06, 
    4.523376e-06, 4.536651e-06, 4.550616e-06, 4.590406e-06, 4.626436e-06, 
    4.665901e-06, 4.675586e-06, 4.722008e-06, 4.684205e-06, 4.746687e-06, 
    4.693545e-06, 4.78575e-06, 4.620801e-06, 4.691978e-06, 4.563474e-06, 
    4.577219e-06, 4.602144e-06, 4.659596e-06, 4.628524e-06, 4.664872e-06, 
    4.584819e-06, 4.543603e-06, 4.532968e-06, 4.513174e-06, 4.533421e-06, 
    4.531772e-06, 4.551192e-06, 4.544946e-06, 4.591731e-06, 4.566566e-06, 
    4.63826e-06, 4.664583e-06, 4.739378e-06, 4.785571e-06, 4.832852e-06, 
    4.853813e-06, 4.860203e-06, 4.862876e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOINTABS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWDP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWLIQ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_DEPTH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SINKS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SOURCES =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1C =
  5.777962, 5.777942, 5.777946, 5.77793, 5.777939, 5.777928, 5.777958, 
    5.777941, 5.777952, 5.77796, 5.777898, 5.777929, 5.777866, 5.777886, 
    5.777836, 5.777869, 5.77783, 5.777837, 5.777814, 5.777821, 5.777792, 
    5.777812, 5.777777, 5.777797, 5.777793, 5.777812, 5.777923, 5.777902, 
    5.777924, 5.777921, 5.777923, 5.777938, 5.777947, 5.777964, 5.777961, 
    5.777948, 5.77792, 5.777929, 5.777905, 5.777905, 5.777878, 5.777891, 
    5.777845, 5.777858, 5.777821, 5.77783, 5.777821, 5.777824, 5.777821, 
    5.777835, 5.777829, 5.777841, 5.777888, 5.777874, 5.777916, 5.777941, 
    5.777957, 5.777969, 5.777967, 5.777965, 5.777948, 5.777933, 5.777921, 
    5.777914, 5.777905, 5.777883, 5.77787, 5.777843, 5.777848, 5.777839, 
    5.777831, 5.777818, 5.77782, 5.777814, 5.777839, 5.777822, 5.77785, 
    5.777843, 5.777904, 5.777927, 5.777936, 5.777945, 5.777966, 5.777952, 
    5.777957, 5.777944, 5.777935, 5.777939, 5.777913, 5.777924, 5.777869, 
    5.777893, 5.777832, 5.777846, 5.777829, 5.777838, 5.777822, 5.777836, 
    5.777812, 5.777806, 5.77781, 5.777796, 5.777837, 5.777821, 5.77794, 
    5.777939, 5.777936, 5.77795, 5.777951, 5.777964, 5.777952, 5.777947, 
    5.777935, 5.777927, 5.77792, 5.777905, 5.777887, 5.777863, 5.777845, 
    5.777834, 5.777841, 5.777835, 5.777842, 5.777845, 5.777808, 5.777829, 
    5.777798, 5.7778, 5.777814, 5.7778, 5.777938, 5.777943, 5.777956, 
    5.777946, 5.777966, 5.777954, 5.777948, 5.777923, 5.777918, 5.777913, 
    5.777903, 5.77789, 5.777868, 5.777848, 5.777831, 5.777832, 5.777832, 
    5.777828, 5.777837, 5.777826, 5.777824, 5.777829, 5.7778, 5.777808, 
    5.7778, 5.777805, 5.777941, 5.777935, 5.777938, 5.777931, 5.777936, 
    5.777915, 5.777908, 5.777878, 5.77789, 5.777871, 5.777888, 5.777885, 
    5.77787, 5.777887, 5.777849, 5.777875, 5.777827, 5.777853, 5.777826, 
    5.777831, 5.777822, 5.777815, 5.777806, 5.777789, 5.777793, 5.777779, 
    5.777925, 5.777915, 5.777916, 5.777907, 5.7779, 5.777886, 5.777862, 
    5.777871, 5.777855, 5.777852, 5.777876, 5.777861, 5.77791, 5.777902, 
    5.777906, 5.777924, 5.777869, 5.777897, 5.777845, 5.777861, 5.777816, 
    5.777838, 5.777795, 5.777776, 5.777759, 5.777739, 5.777911, 5.777917, 
    5.777906, 5.777891, 5.777878, 5.77786, 5.777858, 5.777854, 5.777845, 
    5.777838, 5.777853, 5.777836, 5.7779, 5.777866, 5.777919, 5.777903, 
    5.777892, 5.777897, 5.777872, 5.777866, 5.777842, 5.777854, 5.777781, 
    5.777813, 5.777723, 5.777749, 5.777919, 5.777911, 5.777883, 5.777896, 
    5.777858, 5.777849, 5.777842, 5.777832, 5.777831, 5.777825, 5.777834, 
    5.777825, 5.77786, 5.777844, 5.777886, 5.777876, 5.777881, 5.777886, 
    5.77787, 5.777853, 5.777853, 5.777847, 5.777832, 5.777858, 5.777777, 
    5.777827, 5.777902, 5.777887, 5.777884, 5.777891, 5.77785, 5.777864, 
    5.777825, 5.777836, 5.777818, 5.777827, 5.777828, 5.77784, 5.777846, 
    5.777864, 5.777878, 5.77789, 5.777887, 5.777874, 5.777852, 5.777831, 
    5.777835, 5.77782, 5.777861, 5.777843, 5.777851, 5.777833, 5.777871, 
    5.777839, 5.77788, 5.777876, 5.777865, 5.777843, 5.777838, 5.777833, 
    5.777835, 5.777852, 5.777854, 5.777865, 5.777868, 5.777877, 5.777884, 
    5.777877, 5.777871, 5.777852, 5.777834, 5.777815, 5.777811, 5.777788, 
    5.777806, 5.777777, 5.777802, 5.777758, 5.777837, 5.777802, 5.777864, 
    5.777858, 5.777846, 5.777818, 5.777833, 5.777815, 5.777854, 5.777874, 
    5.777879, 5.777889, 5.777879, 5.77788, 5.77787, 5.777874, 5.777851, 
    5.777863, 5.777828, 5.777816, 5.77778, 5.777758, 5.777736, 5.777726, 
    5.777723, 5.777722 ;

 SOIL1C_TO_SOIL2C =
  3.180418e-08, 3.194395e-08, 3.191678e-08, 3.202952e-08, 3.196698e-08, 
    3.20408e-08, 3.183252e-08, 3.19495e-08, 3.187482e-08, 3.181676e-08, 
    3.224829e-08, 3.203455e-08, 3.24703e-08, 3.233398e-08, 3.267639e-08, 
    3.244909e-08, 3.272223e-08, 3.266983e-08, 3.282751e-08, 3.278234e-08, 
    3.298403e-08, 3.284836e-08, 3.308857e-08, 3.295163e-08, 3.297305e-08, 
    3.284389e-08, 3.207756e-08, 3.222168e-08, 3.206902e-08, 3.208957e-08, 
    3.208035e-08, 3.196827e-08, 3.191179e-08, 3.179349e-08, 3.181497e-08, 
    3.190186e-08, 3.209881e-08, 3.203195e-08, 3.220045e-08, 3.219664e-08, 
    3.238422e-08, 3.229965e-08, 3.261491e-08, 3.252531e-08, 3.278423e-08, 
    3.271911e-08, 3.278117e-08, 3.276235e-08, 3.278141e-08, 3.268592e-08, 
    3.272683e-08, 3.26428e-08, 3.231549e-08, 3.241168e-08, 3.212477e-08, 
    3.195225e-08, 3.183765e-08, 3.175633e-08, 3.176782e-08, 3.178974e-08, 
    3.190236e-08, 3.200825e-08, 3.208894e-08, 3.214291e-08, 3.219609e-08, 
    3.235708e-08, 3.244227e-08, 3.263303e-08, 3.25986e-08, 3.265692e-08, 
    3.271263e-08, 3.280617e-08, 3.279078e-08, 3.283199e-08, 3.265538e-08, 
    3.277276e-08, 3.257899e-08, 3.263199e-08, 3.221056e-08, 3.204999e-08, 
    3.198175e-08, 3.1922e-08, 3.177666e-08, 3.187703e-08, 3.183747e-08, 
    3.19316e-08, 3.199141e-08, 3.196183e-08, 3.214439e-08, 3.207341e-08, 
    3.244732e-08, 3.228627e-08, 3.270614e-08, 3.260567e-08, 3.273022e-08, 
    3.266666e-08, 3.277556e-08, 3.267755e-08, 3.284732e-08, 3.288429e-08, 
    3.285903e-08, 3.295607e-08, 3.267212e-08, 3.278117e-08, 3.196099e-08, 
    3.196582e-08, 3.19883e-08, 3.18895e-08, 3.188345e-08, 3.179291e-08, 
    3.187347e-08, 3.190778e-08, 3.199487e-08, 3.204639e-08, 3.209536e-08, 
    3.220302e-08, 3.232326e-08, 3.24914e-08, 3.261218e-08, 3.269314e-08, 
    3.26435e-08, 3.268733e-08, 3.263833e-08, 3.261536e-08, 3.287044e-08, 
    3.272721e-08, 3.294211e-08, 3.293022e-08, 3.283297e-08, 3.293156e-08, 
    3.196921e-08, 3.194144e-08, 3.184505e-08, 3.192049e-08, 3.178305e-08, 
    3.185998e-08, 3.190422e-08, 3.20749e-08, 3.21124e-08, 3.214717e-08, 
    3.221584e-08, 3.230397e-08, 3.245858e-08, 3.259309e-08, 3.271587e-08, 
    3.270688e-08, 3.271004e-08, 3.273748e-08, 3.266953e-08, 3.274863e-08, 
    3.276191e-08, 3.27272e-08, 3.292863e-08, 3.287108e-08, 3.292997e-08, 
    3.28925e-08, 3.195047e-08, 3.199719e-08, 3.197194e-08, 3.201941e-08, 
    3.198597e-08, 3.213467e-08, 3.217925e-08, 3.238785e-08, 3.230224e-08, 
    3.243849e-08, 3.231608e-08, 3.233777e-08, 3.244294e-08, 3.232269e-08, 
    3.258567e-08, 3.240739e-08, 3.273854e-08, 3.256052e-08, 3.27497e-08, 
    3.271535e-08, 3.277222e-08, 3.282317e-08, 3.288725e-08, 3.300551e-08, 
    3.297812e-08, 3.307701e-08, 3.206683e-08, 3.212742e-08, 3.212208e-08, 
    3.218549e-08, 3.223238e-08, 3.233402e-08, 3.249702e-08, 3.243573e-08, 
    3.254826e-08, 3.257085e-08, 3.239989e-08, 3.250486e-08, 3.216797e-08, 
    3.22224e-08, 3.218999e-08, 3.207161e-08, 3.244985e-08, 3.225574e-08, 
    3.261418e-08, 3.250902e-08, 3.28159e-08, 3.266329e-08, 3.296305e-08, 
    3.30912e-08, 3.321179e-08, 3.335272e-08, 3.216049e-08, 3.211931e-08, 
    3.219303e-08, 3.229502e-08, 3.238964e-08, 3.251544e-08, 3.252831e-08, 
    3.255187e-08, 3.261292e-08, 3.266424e-08, 3.255933e-08, 3.267711e-08, 
    3.223503e-08, 3.24667e-08, 3.210375e-08, 3.221305e-08, 3.228901e-08, 
    3.225568e-08, 3.242872e-08, 3.24695e-08, 3.263522e-08, 3.254956e-08, 
    3.305957e-08, 3.283393e-08, 3.346003e-08, 3.328507e-08, 3.210493e-08, 
    3.216034e-08, 3.235319e-08, 3.226143e-08, 3.252384e-08, 3.258842e-08, 
    3.264093e-08, 3.270804e-08, 3.271529e-08, 3.275505e-08, 3.268989e-08, 
    3.275248e-08, 3.251571e-08, 3.262151e-08, 3.233114e-08, 3.240182e-08, 
    3.236931e-08, 3.233365e-08, 3.244372e-08, 3.256098e-08, 3.256348e-08, 
    3.260108e-08, 3.270705e-08, 3.25249e-08, 3.30887e-08, 3.274052e-08, 
    3.222076e-08, 3.23275e-08, 3.234274e-08, 3.230139e-08, 3.258195e-08, 
    3.248029e-08, 3.275408e-08, 3.268009e-08, 3.280133e-08, 3.274108e-08, 
    3.273222e-08, 3.265484e-08, 3.260667e-08, 3.248496e-08, 3.238592e-08, 
    3.230739e-08, 3.232565e-08, 3.241192e-08, 3.256815e-08, 3.271595e-08, 
    3.268357e-08, 3.279212e-08, 3.250481e-08, 3.262528e-08, 3.257872e-08, 
    3.270013e-08, 3.24341e-08, 3.266065e-08, 3.237619e-08, 3.240113e-08, 
    3.247828e-08, 3.263346e-08, 3.266778e-08, 3.270445e-08, 3.268182e-08, 
    3.257212e-08, 3.255414e-08, 3.24764e-08, 3.245494e-08, 3.23957e-08, 
    3.234666e-08, 3.239147e-08, 3.243852e-08, 3.257216e-08, 3.269259e-08, 
    3.282389e-08, 3.285602e-08, 3.300944e-08, 3.288456e-08, 3.309064e-08, 
    3.291544e-08, 3.321871e-08, 3.267377e-08, 3.291028e-08, 3.248179e-08, 
    3.252795e-08, 3.261145e-08, 3.280295e-08, 3.269956e-08, 3.282047e-08, 
    3.255344e-08, 3.24149e-08, 3.237905e-08, 3.231217e-08, 3.238058e-08, 
    3.237501e-08, 3.244047e-08, 3.241944e-08, 3.25766e-08, 3.249218e-08, 
    3.2732e-08, 3.281951e-08, 3.306665e-08, 3.321815e-08, 3.337236e-08, 
    3.344044e-08, 3.346116e-08, 3.346982e-08 ;

 SOIL1C_TO_SOIL3C =
  3.772076e-10, 3.788659e-10, 3.785436e-10, 3.798811e-10, 3.791391e-10, 
    3.80015e-10, 3.775438e-10, 3.789318e-10, 3.780457e-10, 3.773569e-10, 
    3.824769e-10, 3.799408e-10, 3.851109e-10, 3.834936e-10, 3.875563e-10, 
    3.848593e-10, 3.881002e-10, 3.874785e-10, 3.893494e-10, 3.888135e-10, 
    3.912066e-10, 3.895968e-10, 3.92447e-10, 3.908221e-10, 3.910763e-10, 
    3.895437e-10, 3.804511e-10, 3.821611e-10, 3.803498e-10, 3.805937e-10, 
    3.804842e-10, 3.791545e-10, 3.784844e-10, 3.770808e-10, 3.773356e-10, 
    3.783665e-10, 3.807033e-10, 3.7991e-10, 3.819092e-10, 3.81864e-10, 
    3.840896e-10, 3.830862e-10, 3.868268e-10, 3.857637e-10, 3.888358e-10, 
    3.880632e-10, 3.887995e-10, 3.885763e-10, 3.888024e-10, 3.876693e-10, 
    3.881548e-10, 3.871577e-10, 3.832741e-10, 3.844155e-10, 3.810113e-10, 
    3.789644e-10, 3.776047e-10, 3.766399e-10, 3.767762e-10, 3.770363e-10, 
    3.783725e-10, 3.796288e-10, 3.805861e-10, 3.812266e-10, 3.818575e-10, 
    3.837676e-10, 3.847784e-10, 3.870418e-10, 3.866333e-10, 3.873253e-10, 
    3.879863e-10, 3.890962e-10, 3.889135e-10, 3.894025e-10, 3.87307e-10, 
    3.886997e-10, 3.864006e-10, 3.870295e-10, 3.820292e-10, 3.80124e-10, 
    3.793144e-10, 3.786055e-10, 3.768811e-10, 3.78072e-10, 3.776025e-10, 
    3.787193e-10, 3.79429e-10, 3.79078e-10, 3.812441e-10, 3.80402e-10, 
    3.848383e-10, 3.829275e-10, 3.879093e-10, 3.867171e-10, 3.88195e-10, 
    3.874409e-10, 3.88733e-10, 3.875701e-10, 3.895845e-10, 3.900232e-10, 
    3.897234e-10, 3.908748e-10, 3.875056e-10, 3.887995e-10, 3.790681e-10, 
    3.791254e-10, 3.793921e-10, 3.782198e-10, 3.781481e-10, 3.770738e-10, 
    3.780297e-10, 3.784368e-10, 3.794701e-10, 3.800813e-10, 3.806623e-10, 
    3.819397e-10, 3.833664e-10, 3.853613e-10, 3.867944e-10, 3.877551e-10, 
    3.87166e-10, 3.876861e-10, 3.871047e-10, 3.868322e-10, 3.898588e-10, 
    3.881593e-10, 3.907092e-10, 3.905681e-10, 3.894142e-10, 3.90584e-10, 
    3.791656e-10, 3.788362e-10, 3.776925e-10, 3.785876e-10, 3.769569e-10, 
    3.778697e-10, 3.783945e-10, 3.804196e-10, 3.808645e-10, 3.81277e-10, 
    3.820919e-10, 3.831375e-10, 3.849719e-10, 3.865679e-10, 3.880248e-10, 
    3.879181e-10, 3.879556e-10, 3.882811e-10, 3.874749e-10, 3.884135e-10, 
    3.88571e-10, 3.881591e-10, 3.905492e-10, 3.898664e-10, 3.905651e-10, 
    3.901205e-10, 3.789432e-10, 3.794975e-10, 3.79198e-10, 3.797612e-10, 
    3.793645e-10, 3.811287e-10, 3.816577e-10, 3.841328e-10, 3.83117e-10, 
    3.847336e-10, 3.832812e-10, 3.835385e-10, 3.847864e-10, 3.833596e-10, 
    3.864799e-10, 3.843645e-10, 3.882938e-10, 3.861814e-10, 3.884262e-10, 
    3.880185e-10, 3.886934e-10, 3.892979e-10, 3.900583e-10, 3.914614e-10, 
    3.911365e-10, 3.923099e-10, 3.803238e-10, 3.810427e-10, 3.809794e-10, 
    3.817317e-10, 3.822881e-10, 3.83494e-10, 3.854281e-10, 3.847008e-10, 
    3.86036e-10, 3.86304e-10, 3.842755e-10, 3.85521e-10, 3.815238e-10, 
    3.821697e-10, 3.817851e-10, 3.803805e-10, 3.848684e-10, 3.825653e-10, 
    3.868181e-10, 3.855705e-10, 3.892117e-10, 3.874009e-10, 3.909576e-10, 
    3.924782e-10, 3.939091e-10, 3.955815e-10, 3.81435e-10, 3.809466e-10, 
    3.818212e-10, 3.830313e-10, 3.84154e-10, 3.856466e-10, 3.857993e-10, 
    3.860789e-10, 3.868031e-10, 3.874121e-10, 3.861673e-10, 3.875648e-10, 
    3.823195e-10, 3.850683e-10, 3.807619e-10, 3.820587e-10, 3.829599e-10, 
    3.825646e-10, 3.846176e-10, 3.851015e-10, 3.870679e-10, 3.860514e-10, 
    3.921029e-10, 3.894256e-10, 3.968547e-10, 3.947786e-10, 3.807759e-10, 
    3.814333e-10, 3.837215e-10, 3.826328e-10, 3.857462e-10, 3.865125e-10, 
    3.871355e-10, 3.879319e-10, 3.880178e-10, 3.884897e-10, 3.877165e-10, 
    3.884591e-10, 3.856497e-10, 3.869052e-10, 3.834599e-10, 3.842985e-10, 
    3.839127e-10, 3.834895e-10, 3.847955e-10, 3.861869e-10, 3.862166e-10, 
    3.866628e-10, 3.879201e-10, 3.857588e-10, 3.924486e-10, 3.883173e-10, 
    3.821503e-10, 3.834166e-10, 3.835975e-10, 3.831069e-10, 3.864357e-10, 
    3.852296e-10, 3.884782e-10, 3.876002e-10, 3.890387e-10, 3.883239e-10, 
    3.882187e-10, 3.873006e-10, 3.86729e-10, 3.852849e-10, 3.841099e-10, 
    3.83178e-10, 3.833947e-10, 3.844183e-10, 3.86272e-10, 3.880256e-10, 
    3.876415e-10, 3.889294e-10, 3.855204e-10, 3.869499e-10, 3.863974e-10, 
    3.87838e-10, 3.846815e-10, 3.873696e-10, 3.839944e-10, 3.842903e-10, 
    3.852056e-10, 3.870469e-10, 3.874542e-10, 3.878892e-10, 3.876207e-10, 
    3.863191e-10, 3.861058e-10, 3.851834e-10, 3.849287e-10, 3.842258e-10, 
    3.836439e-10, 3.841756e-10, 3.84734e-10, 3.863196e-10, 3.877486e-10, 
    3.893065e-10, 3.896877e-10, 3.915081e-10, 3.900263e-10, 3.924716e-10, 
    3.903927e-10, 3.939913e-10, 3.875253e-10, 3.903315e-10, 3.852473e-10, 
    3.85795e-10, 3.867857e-10, 3.89058e-10, 3.878312e-10, 3.892659e-10, 
    3.860975e-10, 3.844536e-10, 3.840283e-10, 3.832347e-10, 3.840464e-10, 
    3.839804e-10, 3.847571e-10, 3.845075e-10, 3.863723e-10, 3.853706e-10, 
    3.882161e-10, 3.892545e-10, 3.921869e-10, 3.939846e-10, 3.958144e-10, 
    3.966222e-10, 3.968681e-10, 3.969709e-10 ;

 SOIL1C_vr =
  19.97934, 19.97928, 19.97929, 19.97925, 19.97927, 19.97925, 19.97933, 
    19.97928, 19.97931, 19.97933, 19.97917, 19.97925, 19.97908, 19.97913, 
    19.979, 19.97909, 19.97898, 19.979, 19.97894, 19.97896, 19.97888, 
    19.97894, 19.97884, 19.9789, 19.97889, 19.97894, 19.97923, 19.97918, 
    19.97923, 19.97923, 19.97923, 19.97927, 19.9793, 19.97934, 19.97933, 
    19.9793, 19.97922, 19.97925, 19.97918, 19.97919, 19.97911, 19.97915, 
    19.97902, 19.97906, 19.97896, 19.97898, 19.97896, 19.97897, 19.97896, 
    19.979, 19.97898, 19.97901, 19.97914, 19.9791, 19.97921, 19.97928, 
    19.97932, 19.97935, 19.97935, 19.97934, 19.9793, 19.97926, 19.97923, 
    19.97921, 19.97919, 19.97912, 19.97909, 19.97902, 19.97903, 19.97901, 
    19.97899, 19.97895, 19.97896, 19.97894, 19.97901, 19.97896, 19.97904, 
    19.97902, 19.97918, 19.97924, 19.97927, 19.97929, 19.97935, 19.97931, 
    19.97932, 19.97929, 19.97927, 19.97928, 19.97921, 19.97923, 19.97909, 
    19.97915, 19.97899, 19.97903, 19.97898, 19.979, 19.97896, 19.979, 
    19.97894, 19.97892, 19.97893, 19.97889, 19.979, 19.97896, 19.97928, 
    19.97927, 19.97927, 19.9793, 19.97931, 19.97934, 19.97931, 19.9793, 
    19.97926, 19.97924, 19.97923, 19.97918, 19.97914, 19.97907, 19.97902, 
    19.97899, 19.97901, 19.979, 19.97902, 19.97902, 19.97893, 19.97898, 
    19.9789, 19.9789, 19.97894, 19.9789, 19.97927, 19.97928, 19.97932, 
    19.97929, 19.97935, 19.97931, 19.9793, 19.97923, 19.97922, 19.9792, 
    19.97918, 19.97914, 19.97908, 19.97903, 19.97898, 19.97899, 19.97899, 
    19.97898, 19.979, 19.97897, 19.97897, 19.97898, 19.9789, 19.97893, 
    19.9789, 19.97892, 19.97928, 19.97926, 19.97927, 19.97925, 19.97927, 
    19.97921, 19.97919, 19.97911, 19.97915, 19.97909, 19.97914, 19.97913, 
    19.97909, 19.97914, 19.97904, 19.9791, 19.97898, 19.97905, 19.97897, 
    19.97899, 19.97896, 19.97894, 19.97892, 19.97887, 19.97889, 19.97885, 
    19.97923, 19.97921, 19.97921, 19.97919, 19.97917, 19.97913, 19.97907, 
    19.97909, 19.97905, 19.97904, 19.97911, 19.97907, 19.9792, 19.97918, 
    19.97919, 19.97923, 19.97909, 19.97916, 19.97902, 19.97906, 19.97895, 
    19.97901, 19.97889, 19.97884, 19.9788, 19.97874, 19.9792, 19.97922, 
    19.97919, 19.97915, 19.97911, 19.97906, 19.97906, 19.97905, 19.97902, 
    19.97901, 19.97905, 19.979, 19.97917, 19.97908, 19.97922, 19.97918, 
    19.97915, 19.97916, 19.9791, 19.97908, 19.97902, 19.97905, 19.97885, 
    19.97894, 19.9787, 19.97877, 19.97922, 19.9792, 19.97912, 19.97916, 
    19.97906, 19.97903, 19.97902, 19.97899, 19.97899, 19.97897, 19.979, 
    19.97897, 19.97906, 19.97902, 19.97913, 19.97911, 19.97912, 19.97913, 
    19.97909, 19.97905, 19.97904, 19.97903, 19.97899, 19.97906, 19.97884, 
    19.97898, 19.97918, 19.97914, 19.97913, 19.97915, 19.97904, 19.97908, 
    19.97897, 19.979, 19.97895, 19.97898, 19.97898, 19.97901, 19.97903, 
    19.97907, 19.97911, 19.97914, 19.97914, 19.9791, 19.97904, 19.97898, 
    19.979, 19.97896, 19.97907, 19.97902, 19.97904, 19.97899, 19.97909, 
    19.97901, 19.97912, 19.97911, 19.97908, 19.97902, 19.979, 19.97899, 
    19.979, 19.97904, 19.97905, 19.97908, 19.97909, 19.97911, 19.97913, 
    19.97911, 19.97909, 19.97904, 19.97899, 19.97894, 19.97893, 19.97887, 
    19.97892, 19.97884, 19.97891, 19.97879, 19.979, 19.97891, 19.97908, 
    19.97906, 19.97902, 19.97895, 19.97899, 19.97894, 19.97905, 19.9791, 
    19.97911, 19.97914, 19.97911, 19.97912, 19.97909, 19.9791, 19.97904, 
    19.97907, 19.97898, 19.97895, 19.97885, 19.97879, 19.97873, 19.97871, 
    19.9787, 19.9787,
  19.981, 19.98093, 19.98095, 19.98089, 19.98092, 19.98088, 19.98099, 
    19.98093, 19.98097, 19.981, 19.98078, 19.98089, 19.98067, 19.98074, 
    19.98056, 19.98068, 19.98054, 19.98057, 19.98049, 19.98051, 19.98041, 
    19.98048, 19.98036, 19.98042, 19.98041, 19.98048, 19.98087, 19.98079, 
    19.98087, 19.98086, 19.98087, 19.98092, 19.98095, 19.98101, 19.981, 
    19.98096, 19.98086, 19.98089, 19.9808, 19.98081, 19.98071, 19.98075, 
    19.98059, 19.98064, 19.98051, 19.98054, 19.98051, 19.98052, 19.98051, 
    19.98056, 19.98054, 19.98058, 19.98075, 19.9807, 19.98084, 19.98093, 
    19.98099, 19.98103, 19.98102, 19.98101, 19.98096, 19.9809, 19.98086, 
    19.98083, 19.98081, 19.98072, 19.98068, 19.98059, 19.9806, 19.98057, 
    19.98055, 19.9805, 19.9805, 19.98048, 19.98057, 19.98051, 19.98061, 
    19.98059, 19.9808, 19.98088, 19.98092, 19.98095, 19.98102, 19.98097, 
    19.98099, 19.98094, 19.98091, 19.98092, 19.98083, 19.98087, 19.98068, 
    19.98076, 19.98055, 19.9806, 19.98054, 19.98057, 19.98051, 19.98056, 
    19.98048, 19.98046, 19.98047, 19.98042, 19.98057, 19.98051, 19.98093, 
    19.98092, 19.98091, 19.98096, 19.98096, 19.98101, 19.98097, 19.98095, 
    19.98091, 19.98088, 19.98086, 19.9808, 19.98074, 19.98066, 19.9806, 
    19.98055, 19.98058, 19.98056, 19.98058, 19.98059, 19.98046, 19.98054, 
    19.98043, 19.98043, 19.98048, 19.98043, 19.98092, 19.98094, 19.98099, 
    19.98095, 19.98102, 19.98098, 19.98096, 19.98087, 19.98085, 19.98083, 
    19.9808, 19.98075, 19.98067, 19.98061, 19.98054, 19.98055, 19.98055, 
    19.98053, 19.98057, 19.98053, 19.98052, 19.98054, 19.98044, 19.98046, 
    19.98043, 19.98045, 19.98093, 19.98091, 19.98092, 19.9809, 19.98091, 
    19.98084, 19.98082, 19.98071, 19.98075, 19.98068, 19.98075, 19.98073, 
    19.98068, 19.98074, 19.98061, 19.9807, 19.98053, 19.98062, 19.98053, 
    19.98054, 19.98051, 19.98049, 19.98046, 19.9804, 19.98041, 19.98036, 
    19.98087, 19.98084, 19.98084, 19.98081, 19.98079, 19.98074, 19.98065, 
    19.98068, 19.98063, 19.98062, 19.9807, 19.98065, 19.98082, 19.98079, 
    19.98081, 19.98087, 19.98068, 19.98078, 19.98059, 19.98065, 19.98049, 
    19.98057, 19.98042, 19.98035, 19.98029, 19.98022, 19.98083, 19.98084, 
    19.98081, 19.98076, 19.98071, 19.98064, 19.98064, 19.98063, 19.98059, 
    19.98057, 19.98062, 19.98056, 19.98079, 19.98067, 19.98085, 19.9808, 
    19.98076, 19.98078, 19.98069, 19.98067, 19.98058, 19.98063, 19.98037, 
    19.98048, 19.98017, 19.98026, 19.98085, 19.98083, 19.98073, 19.98077, 
    19.98064, 19.98061, 19.98058, 19.98055, 19.98054, 19.98052, 19.98056, 
    19.98052, 19.98064, 19.98059, 19.98074, 19.9807, 19.98072, 19.98074, 
    19.98068, 19.98062, 19.98062, 19.9806, 19.98055, 19.98064, 19.98036, 
    19.98053, 19.98079, 19.98074, 19.98073, 19.98075, 19.98061, 19.98066, 
    19.98052, 19.98056, 19.9805, 19.98053, 19.98054, 19.98057, 19.9806, 
    19.98066, 19.98071, 19.98075, 19.98074, 19.9807, 19.98062, 19.98054, 
    19.98056, 19.9805, 19.98065, 19.98059, 19.98061, 19.98055, 19.98069, 
    19.98057, 19.98071, 19.9807, 19.98066, 19.98059, 19.98057, 19.98055, 
    19.98056, 19.98062, 19.98063, 19.98067, 19.98067, 19.98071, 19.98073, 
    19.98071, 19.98068, 19.98062, 19.98055, 19.98049, 19.98047, 19.98039, 
    19.98046, 19.98035, 19.98044, 19.98029, 19.98056, 19.98045, 19.98066, 
    19.98064, 19.9806, 19.9805, 19.98055, 19.98049, 19.98063, 19.9807, 
    19.98071, 19.98075, 19.98071, 19.98072, 19.98068, 19.98069, 19.98061, 
    19.98066, 19.98054, 19.98049, 19.98037, 19.98029, 19.98021, 19.98018, 
    19.98017, 19.98016,
  19.98273, 19.98265, 19.98267, 19.9826, 19.98264, 19.9826, 19.98271, 
    19.98265, 19.98269, 19.98272, 19.98249, 19.9826, 19.98237, 19.98244, 
    19.98226, 19.98238, 19.98223, 19.98226, 19.98217, 19.9822, 19.98209, 
    19.98216, 19.98203, 19.98211, 19.9821, 19.98217, 19.98258, 19.9825, 
    19.98258, 19.98257, 19.98258, 19.98264, 19.98267, 19.98273, 19.98272, 
    19.98268, 19.98257, 19.9826, 19.98251, 19.98252, 19.98241, 19.98246, 
    19.98229, 19.98234, 19.9822, 19.98223, 19.9822, 19.98221, 19.9822, 
    19.98225, 19.98223, 19.98228, 19.98245, 19.9824, 19.98255, 19.98265, 
    19.98271, 19.98275, 19.98275, 19.98274, 19.98268, 19.98262, 19.98257, 
    19.98254, 19.98252, 19.98243, 19.98238, 19.98228, 19.9823, 19.98227, 
    19.98224, 19.98219, 19.98219, 19.98217, 19.98227, 19.9822, 19.98231, 
    19.98228, 19.98251, 19.9826, 19.98263, 19.98266, 19.98274, 19.98269, 
    19.98271, 19.98266, 19.98263, 19.98264, 19.98254, 19.98258, 19.98238, 
    19.98247, 19.98224, 19.98229, 19.98223, 19.98226, 19.9822, 19.98226, 
    19.98216, 19.98214, 19.98216, 19.98211, 19.98226, 19.9822, 19.98264, 
    19.98264, 19.98263, 19.98268, 19.98269, 19.98273, 19.98269, 19.98267, 
    19.98262, 19.9826, 19.98257, 19.98251, 19.98245, 19.98236, 19.98229, 
    19.98225, 19.98227, 19.98225, 19.98228, 19.98229, 19.98215, 19.98223, 
    19.98211, 19.98212, 19.98217, 19.98212, 19.98264, 19.98265, 19.98271, 
    19.98266, 19.98274, 19.9827, 19.98267, 19.98258, 19.98256, 19.98254, 
    19.98251, 19.98246, 19.98237, 19.9823, 19.98223, 19.98224, 19.98224, 
    19.98222, 19.98226, 19.98222, 19.98221, 19.98223, 19.98212, 19.98215, 
    19.98212, 19.98214, 19.98265, 19.98262, 19.98264, 19.98261, 19.98263, 
    19.98255, 19.98252, 19.98241, 19.98246, 19.98238, 19.98245, 19.98244, 
    19.98238, 19.98245, 19.98231, 19.9824, 19.98222, 19.98232, 19.98222, 
    19.98223, 19.9822, 19.98218, 19.98214, 19.98208, 19.98209, 19.98204, 
    19.98259, 19.98255, 19.98256, 19.98252, 19.9825, 19.98244, 19.98235, 
    19.98239, 19.98232, 19.98231, 19.9824, 19.98235, 19.98253, 19.9825, 
    19.98252, 19.98258, 19.98238, 19.98248, 19.98229, 19.98235, 19.98218, 
    19.98226, 19.9821, 19.98203, 19.98197, 19.98189, 19.98253, 19.98256, 
    19.98252, 19.98246, 19.98241, 19.98234, 19.98234, 19.98232, 19.98229, 
    19.98226, 19.98232, 19.98226, 19.98249, 19.98237, 19.98256, 19.98251, 
    19.98247, 19.98248, 19.98239, 19.98237, 19.98228, 19.98232, 19.98205, 
    19.98217, 19.98183, 19.98193, 19.98256, 19.98253, 19.98243, 19.98248, 
    19.98234, 19.9823, 19.98228, 19.98224, 19.98223, 19.98221, 19.98225, 
    19.98221, 19.98234, 19.98229, 19.98244, 19.9824, 19.98242, 19.98244, 
    19.98238, 19.98232, 19.98232, 19.9823, 19.98224, 19.98234, 19.98203, 
    19.98222, 19.9825, 19.98244, 19.98244, 19.98246, 19.98231, 19.98236, 
    19.98221, 19.98225, 19.98219, 19.98222, 19.98223, 19.98227, 19.98229, 
    19.98236, 19.98241, 19.98246, 19.98244, 19.9824, 19.98232, 19.98223, 
    19.98225, 19.98219, 19.98235, 19.98228, 19.98231, 19.98224, 19.98239, 
    19.98226, 19.98242, 19.9824, 19.98236, 19.98228, 19.98226, 19.98224, 
    19.98225, 19.98231, 19.98232, 19.98236, 19.98238, 19.98241, 19.98243, 
    19.98241, 19.98238, 19.98231, 19.98225, 19.98218, 19.98216, 19.98208, 
    19.98214, 19.98203, 19.98213, 19.98196, 19.98226, 19.98213, 19.98236, 
    19.98234, 19.98229, 19.98219, 19.98224, 19.98218, 19.98232, 19.9824, 
    19.98242, 19.98245, 19.98242, 19.98242, 19.98238, 19.9824, 19.98231, 
    19.98236, 19.98223, 19.98218, 19.98205, 19.98196, 19.98188, 19.98184, 
    19.98183, 19.98183,
  19.9841, 19.98403, 19.98404, 19.98398, 19.98401, 19.98397, 19.98409, 
    19.98402, 19.98406, 19.98409, 19.98386, 19.98398, 19.98375, 19.98382, 
    19.98363, 19.98376, 19.98361, 19.98364, 19.98355, 19.98358, 19.98347, 
    19.98354, 19.98341, 19.98349, 19.98347, 19.98355, 19.98396, 19.98388, 
    19.98396, 19.98395, 19.98395, 19.98401, 19.98405, 19.98411, 19.9841, 
    19.98405, 19.98394, 19.98398, 19.98389, 19.98389, 19.98379, 19.98384, 
    19.98367, 19.98372, 19.98358, 19.98361, 19.98358, 19.98359, 19.98358, 
    19.98363, 19.98361, 19.98365, 19.98383, 19.98378, 19.98393, 19.98402, 
    19.98409, 19.98413, 19.98412, 19.98411, 19.98405, 19.98399, 19.98395, 
    19.98392, 19.98389, 19.9838, 19.98376, 19.98366, 19.98368, 19.98364, 
    19.98361, 19.98356, 19.98357, 19.98355, 19.98365, 19.98358, 19.98369, 
    19.98366, 19.98388, 19.98397, 19.98401, 19.98404, 19.98412, 19.98406, 
    19.98409, 19.98403, 19.984, 19.98402, 19.98392, 19.98396, 19.98376, 
    19.98384, 19.98362, 19.98367, 19.98361, 19.98364, 19.98358, 19.98363, 
    19.98354, 19.98352, 19.98354, 19.98348, 19.98364, 19.98358, 19.98402, 
    19.98402, 19.984, 19.98406, 19.98406, 19.98411, 19.98407, 19.98405, 
    19.984, 19.98397, 19.98395, 19.98389, 19.98382, 19.98373, 19.98367, 
    19.98363, 19.98365, 19.98363, 19.98365, 19.98367, 19.98353, 19.98361, 
    19.98349, 19.9835, 19.98355, 19.9835, 19.98401, 19.98403, 19.98408, 
    19.98404, 19.98411, 19.98407, 19.98405, 19.98396, 19.98394, 19.98392, 
    19.98388, 19.98383, 19.98375, 19.98368, 19.98361, 19.98362, 19.98362, 
    19.9836, 19.98364, 19.98359, 19.98359, 19.98361, 19.9835, 19.98353, 
    19.9835, 19.98352, 19.98402, 19.984, 19.98401, 19.98399, 19.984, 
    19.98392, 19.9839, 19.98379, 19.98384, 19.98376, 19.98383, 19.98382, 
    19.98376, 19.98382, 19.98368, 19.98378, 19.9836, 19.9837, 19.98359, 
    19.98361, 19.98358, 19.98355, 19.98352, 19.98346, 19.98347, 19.98342, 
    19.98396, 19.98393, 19.98393, 19.9839, 19.98387, 19.98382, 19.98373, 
    19.98376, 19.9837, 19.98369, 19.98378, 19.98373, 19.98391, 19.98388, 
    19.98389, 19.98396, 19.98376, 19.98386, 19.98367, 19.98372, 19.98356, 
    19.98364, 19.98348, 19.98341, 19.98335, 19.98327, 19.98391, 19.98393, 
    19.98389, 19.98384, 19.98379, 19.98372, 19.98371, 19.9837, 19.98367, 
    19.98364, 19.9837, 19.98363, 19.98387, 19.98375, 19.98394, 19.98388, 
    19.98384, 19.98386, 19.98377, 19.98375, 19.98366, 19.9837, 19.98343, 
    19.98355, 19.98322, 19.98331, 19.98394, 19.98391, 19.98381, 19.98386, 
    19.98372, 19.98368, 19.98365, 19.98362, 19.98361, 19.98359, 19.98363, 
    19.98359, 19.98372, 19.98366, 19.98382, 19.98378, 19.9838, 19.98382, 
    19.98376, 19.9837, 19.98369, 19.98368, 19.98362, 19.98372, 19.98341, 
    19.9836, 19.98388, 19.98382, 19.98381, 19.98384, 19.98368, 19.98374, 
    19.98359, 19.98363, 19.98357, 19.9836, 19.9836, 19.98365, 19.98367, 
    19.98374, 19.98379, 19.98383, 19.98382, 19.98378, 19.98369, 19.98361, 
    19.98363, 19.98357, 19.98373, 19.98366, 19.98369, 19.98362, 19.98376, 
    19.98364, 19.9838, 19.98378, 19.98374, 19.98366, 19.98364, 19.98362, 
    19.98363, 19.98369, 19.9837, 19.98374, 19.98375, 19.98379, 19.98381, 
    19.98379, 19.98376, 19.98369, 19.98363, 19.98355, 19.98354, 19.98346, 
    19.98352, 19.98341, 19.98351, 19.98334, 19.98363, 19.98351, 19.98374, 
    19.98371, 19.98367, 19.98357, 19.98362, 19.98356, 19.9837, 19.98377, 
    19.98379, 19.98383, 19.98379, 19.9838, 19.98376, 19.98377, 19.98369, 
    19.98373, 19.9836, 19.98356, 19.98343, 19.98334, 19.98326, 19.98322, 
    19.98321, 19.98321,
  19.98571, 19.98564, 19.98565, 19.9856, 19.98563, 19.98559, 19.98569, 
    19.98564, 19.98567, 19.9857, 19.98549, 19.9856, 19.98539, 19.98545, 
    19.98529, 19.9854, 19.98527, 19.98529, 19.98522, 19.98524, 19.98514, 
    19.98521, 19.98509, 19.98516, 19.98515, 19.98521, 19.98558, 19.98551, 
    19.98558, 19.98557, 19.98557, 19.98563, 19.98565, 19.98571, 19.9857, 
    19.98566, 19.98557, 19.9856, 19.98552, 19.98552, 19.98543, 19.98547, 
    19.98532, 19.98536, 19.98524, 19.98527, 19.98524, 19.98525, 19.98524, 
    19.98529, 19.98527, 19.98531, 19.98546, 19.98542, 19.98555, 19.98564, 
    19.98569, 19.98573, 19.98572, 19.98571, 19.98566, 19.98561, 19.98557, 
    19.98554, 19.98552, 19.98544, 19.9854, 19.98531, 19.98533, 19.9853, 
    19.98527, 19.98523, 19.98524, 19.98522, 19.9853, 19.98524, 19.98534, 
    19.98531, 19.98551, 19.98559, 19.98562, 19.98565, 19.98572, 19.98567, 
    19.98569, 19.98565, 19.98562, 19.98563, 19.98554, 19.98558, 19.9854, 
    19.98548, 19.98528, 19.98532, 19.98527, 19.98529, 19.98524, 19.98529, 
    19.98521, 19.98519, 19.9852, 19.98516, 19.98529, 19.98524, 19.98563, 
    19.98563, 19.98562, 19.98567, 19.98567, 19.98571, 19.98567, 19.98566, 
    19.98561, 19.98559, 19.98557, 19.98552, 19.98546, 19.98538, 19.98532, 
    19.98528, 19.98531, 19.98528, 19.98531, 19.98532, 19.9852, 19.98527, 
    19.98516, 19.98517, 19.98522, 19.98517, 19.98563, 19.98564, 19.98569, 
    19.98565, 19.98572, 19.98568, 19.98566, 19.98558, 19.98556, 19.98554, 
    19.98551, 19.98547, 19.98539, 19.98533, 19.98527, 19.98528, 19.98528, 
    19.98526, 19.98529, 19.98526, 19.98525, 19.98527, 19.98517, 19.9852, 
    19.98517, 19.98519, 19.98564, 19.98561, 19.98563, 19.9856, 19.98562, 
    19.98555, 19.98553, 19.98543, 19.98547, 19.9854, 19.98546, 19.98545, 
    19.9854, 19.98546, 19.98533, 19.98542, 19.98526, 19.98535, 19.98526, 
    19.98527, 19.98524, 19.98522, 19.98519, 19.98513, 19.98515, 19.9851, 
    19.98558, 19.98555, 19.98556, 19.98553, 19.9855, 19.98545, 19.98538, 
    19.9854, 19.98535, 19.98534, 19.98542, 19.98537, 19.98553, 19.98551, 
    19.98552, 19.98558, 19.9854, 19.98549, 19.98532, 19.98537, 19.98522, 
    19.9853, 19.98515, 19.98509, 19.98503, 19.98497, 19.98554, 19.98556, 
    19.98552, 19.98547, 19.98543, 19.98537, 19.98536, 19.98535, 19.98532, 
    19.9853, 19.98535, 19.98529, 19.9855, 19.98539, 19.98556, 19.98551, 
    19.98548, 19.98549, 19.98541, 19.98539, 19.98531, 19.98535, 19.98511, 
    19.98522, 19.98492, 19.985, 19.98556, 19.98554, 19.98545, 19.98549, 
    19.98536, 19.98533, 19.98531, 19.98528, 19.98527, 19.98525, 19.98528, 
    19.98525, 19.98537, 19.98532, 19.98545, 19.98542, 19.98544, 19.98545, 
    19.9854, 19.98535, 19.98534, 19.98533, 19.98528, 19.98536, 19.98509, 
    19.98526, 19.98551, 19.98546, 19.98545, 19.98547, 19.98534, 19.98538, 
    19.98525, 19.98529, 19.98523, 19.98526, 19.98526, 19.9853, 19.98532, 
    19.98538, 19.98543, 19.98547, 19.98546, 19.98542, 19.98534, 19.98527, 
    19.98529, 19.98524, 19.98537, 19.98532, 19.98534, 19.98528, 19.98541, 
    19.9853, 19.98543, 19.98542, 19.98539, 19.98531, 19.98529, 19.98528, 
    19.98529, 19.98534, 19.98535, 19.98539, 19.9854, 19.98542, 19.98545, 
    19.98543, 19.9854, 19.98534, 19.98528, 19.98522, 19.9852, 19.98513, 
    19.98519, 19.98509, 19.98518, 19.98503, 19.98529, 19.98518, 19.98538, 
    19.98536, 19.98532, 19.98523, 19.98528, 19.98522, 19.98535, 19.98541, 
    19.98543, 19.98546, 19.98543, 19.98543, 19.9854, 19.98541, 19.98534, 
    19.98538, 19.98526, 19.98522, 19.9851, 19.98503, 19.98496, 19.98493, 
    19.98491, 19.98491,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N =
  0.7222453, 0.7222428, 0.7222432, 0.7222412, 0.7222424, 0.722241, 0.7222448, 
    0.7222427, 0.722244, 0.722245, 0.7222373, 0.7222411, 0.7222332, 
    0.7222357, 0.7222295, 0.7222337, 0.7222287, 0.7222297, 0.7222268, 
    0.7222276, 0.722224, 0.7222264, 0.7222221, 0.7222246, 0.7222242, 
    0.7222265, 0.7222403, 0.7222378, 0.7222405, 0.7222401, 0.7222403, 
    0.7222423, 0.7222434, 0.7222455, 0.7222451, 0.7222435, 0.72224, 
    0.7222412, 0.7222381, 0.7222382, 0.7222348, 0.7222363, 0.7222307, 
    0.7222323, 0.7222276, 0.7222288, 0.7222276, 0.722228, 0.7222276, 
    0.7222294, 0.7222286, 0.7222301, 0.722236, 0.7222343, 0.7222395, 
    0.7222426, 0.7222447, 0.7222462, 0.7222459, 0.7222456, 0.7222435, 
    0.7222416, 0.7222401, 0.7222392, 0.7222382, 0.7222353, 0.7222338, 
    0.7222303, 0.722231, 0.7222299, 0.7222289, 0.7222272, 0.7222275, 
    0.7222267, 0.7222299, 0.7222278, 0.7222313, 0.7222303, 0.7222379, 
    0.7222409, 0.7222421, 0.7222431, 0.7222458, 0.722244, 0.7222447, 
    0.722243, 0.7222419, 0.7222424, 0.7222391, 0.7222404, 0.7222337, 
    0.7222366, 0.722229, 0.7222308, 0.7222286, 0.7222297, 0.7222278, 
    0.7222295, 0.7222264, 0.7222258, 0.7222263, 0.7222245, 0.7222296, 
    0.7222276, 0.7222425, 0.7222424, 0.7222419, 0.7222437, 0.7222438, 
    0.7222455, 0.722244, 0.7222434, 0.7222418, 0.7222409, 0.72224, 0.7222381, 
    0.7222359, 0.7222329, 0.7222307, 0.7222292, 0.7222301, 0.7222294, 
    0.7222303, 0.7222306, 0.722226, 0.7222286, 0.7222248, 0.722225, 
    0.7222267, 0.722225, 0.7222423, 0.7222428, 0.7222446, 0.7222432, 
    0.7222457, 0.7222443, 0.7222435, 0.7222404, 0.7222397, 0.7222391, 
    0.7222378, 0.7222363, 0.7222335, 0.722231, 0.7222288, 0.722229, 
    0.7222289, 0.7222285, 0.7222297, 0.7222282, 0.722228, 0.7222286, 
    0.722225, 0.722226, 0.722225, 0.7222257, 0.7222427, 0.7222418, 0.7222422, 
    0.7222414, 0.722242, 0.7222393, 0.7222385, 0.7222347, 0.7222363, 
    0.7222338, 0.722236, 0.7222357, 0.7222338, 0.7222359, 0.7222311, 
    0.7222344, 0.7222284, 0.7222316, 0.7222282, 0.7222288, 0.7222278, 
    0.7222269, 0.7222257, 0.7222236, 0.7222241, 0.7222223, 0.7222406, 
    0.7222394, 0.7222396, 0.7222384, 0.7222375, 0.7222357, 0.7222328, 
    0.7222339, 0.7222319, 0.7222314, 0.7222345, 0.7222326, 0.7222387, 
    0.7222377, 0.7222383, 0.7222404, 0.7222337, 0.7222371, 0.7222307, 
    0.7222326, 0.722227, 0.7222298, 0.7222244, 0.722222, 0.7222199, 
    0.7222173, 0.7222388, 0.7222396, 0.7222382, 0.7222364, 0.7222347, 
    0.7222325, 0.7222322, 0.7222318, 0.7222307, 0.7222298, 0.7222316, 
    0.7222295, 0.7222375, 0.7222333, 0.7222399, 0.7222379, 0.7222365, 
    0.7222371, 0.722234, 0.7222333, 0.7222303, 0.7222318, 0.7222226, 
    0.7222267, 0.7222154, 0.7222186, 0.7222399, 0.7222388, 0.7222354, 
    0.7222371, 0.7222323, 0.7222311, 0.7222302, 0.7222289, 0.7222288, 
    0.7222281, 0.7222293, 0.7222282, 0.7222325, 0.7222306, 0.7222358, 
    0.7222345, 0.7222351, 0.7222357, 0.7222337, 0.7222316, 0.7222316, 
    0.7222309, 0.722229, 0.7222323, 0.7222221, 0.7222284, 0.7222378, 
    0.7222359, 0.7222356, 0.7222363, 0.7222313, 0.7222331, 0.7222281, 
    0.7222295, 0.7222273, 0.7222283, 0.7222285, 0.72223, 0.7222308, 0.722233, 
    0.7222348, 0.7222362, 0.7222359, 0.7222343, 0.7222315, 0.7222288, 
    0.7222294, 0.7222275, 0.7222326, 0.7222304, 0.7222313, 0.7222291, 
    0.7222339, 0.7222298, 0.722235, 0.7222345, 0.7222331, 0.7222303, 
    0.7222297, 0.7222291, 0.7222294, 0.7222314, 0.7222317, 0.7222332, 
    0.7222335, 0.7222346, 0.7222355, 0.7222347, 0.7222338, 0.7222314, 
    0.7222292, 0.7222269, 0.7222263, 0.7222235, 0.7222258, 0.7222221, 
    0.7222252, 0.7222198, 0.7222296, 0.7222253, 0.7222331, 0.7222322, 
    0.7222307, 0.7222273, 0.7222291, 0.7222269, 0.7222317, 0.7222342, 
    0.7222349, 0.7222361, 0.7222349, 0.722235, 0.7222338, 0.7222342, 
    0.7222313, 0.7222329, 0.7222285, 0.722227, 0.7222225, 0.7222198, 
    0.722217, 0.7222158, 0.7222154, 0.7222152 ;

 SOIL1N_TNDNCY_VERT_TRANS =
  -1.027984e-20, 5.139921e-21, -3.597945e-20, -2.569961e-20, 2.006177e-36, 
    -5.139921e-21, 5.139921e-21, 1.027984e-20, 3.083953e-20, -1.541976e-20, 
    -2.055969e-20, 2.055969e-20, -5.139921e-21, 5.139921e-21, -1.027984e-20, 
    5.139921e-21, 0, -1.027984e-20, 1.027984e-20, -1.027984e-20, 
    2.055969e-20, -2.006177e-36, -1.027984e-20, -1.027984e-20, 2.569961e-20, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, 1.027984e-20, -5.139921e-21, 
    -1.541976e-20, 5.139921e-21, -2.055969e-20, -4.111937e-20, -5.139921e-21, 
    1.027984e-20, 0, -1.027984e-20, 2.055969e-20, -1.027984e-20, 
    -2.055969e-20, 2.006177e-36, 0, -3.597945e-20, 1.541976e-20, 
    5.139921e-21, -1.027984e-20, 0, 0, 2.055969e-20, 1.027984e-20, 
    -6.167906e-20, 5.139921e-21, 1.027984e-20, 2.055969e-20, -1.027984e-20, 
    1.027984e-20, -1.027984e-20, -2.055969e-20, -1.541976e-20, -1.027984e-20, 
    -1.027984e-20, 5.139921e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -5.139921e-21, -2.055969e-20, -2.569961e-20, 5.139921e-21, -2.055969e-20, 
    1.027984e-20, 3.083953e-20, -1.541976e-20, 1.027984e-20, 3.083953e-20, 
    2.569961e-20, -1.027984e-20, -4.625929e-20, -3.083953e-20, -1.027984e-20, 
    -1.027984e-20, 5.139921e-21, 1.027984e-20, 2.569961e-20, -1.541976e-20, 
    -5.139921e-21, -1.027984e-20, 0, -1.541976e-20, -2.569961e-20, 
    2.055969e-20, 2.569961e-20, 1.027984e-20, 5.139921e-21, -5.139921e-21, 0, 
    -1.541976e-20, -2.006177e-36, 1.027984e-20, 3.597945e-20, -5.139921e-21, 
    -5.139921e-21, 1.027984e-20, -2.569961e-20, -1.027984e-20, -1.027984e-20, 
    1.541976e-20, -4.111937e-20, 1.541976e-20, 1.027984e-20, -3.597945e-20, 
    -1.027984e-20, 2.055969e-20, -3.597945e-20, -1.541976e-20, 2.055969e-20, 
    1.541976e-20, 2.569961e-20, -5.139921e-21, 4.111937e-20, -1.027984e-20, 
    1.541976e-20, 0, 0, 0, -2.006177e-36, -1.027984e-20, 0, 5.139921e-21, 
    2.055969e-20, -2.569961e-20, -3.083953e-20, 1.027984e-20, 1.541976e-20, 
    -1.541976e-20, 5.139921e-21, -1.541976e-20, 0, 2.569961e-20, 
    -2.055969e-20, -2.055969e-20, -1.027984e-20, 3.083953e-20, -1.541976e-20, 
    -2.569961e-20, 1.541976e-20, 1.027984e-20, -1.027984e-20, -1.027984e-20, 
    5.139921e-21, 5.139921e-21, -5.139921e-21, 0, 0, 2.055969e-20, 
    3.083953e-20, 5.139921e-21, -1.541976e-20, -1.027984e-20, 1.541976e-20, 
    -3.083953e-20, 5.139921e-21, 1.541976e-20, -1.541976e-20, 2.006177e-36, 
    -1.541976e-20, -5.139921e-21, -5.139921e-21, 2.569961e-20, 2.055969e-20, 
    5.139921e-21, -1.541976e-20, 0, -1.541976e-20, 1.027984e-20, 
    -2.055969e-20, 0, -2.006177e-36, -5.139921e-21, 1.027984e-20, 
    2.569961e-20, 3.083953e-20, -5.139921e-21, -1.027984e-20, 5.139921e-21, 
    1.027984e-20, 5.139921e-21, 1.027984e-20, 5.139921e-21, -1.541976e-20, 
    2.006177e-36, -1.027984e-20, 5.139921e-21, 5.139921e-21, -2.569961e-20, 
    5.139921e-21, 1.541976e-20, -1.541976e-20, -1.541976e-20, 0, 
    -3.597945e-20, 1.027984e-20, -1.541976e-20, -1.027984e-20, 2.055969e-20, 
    2.055969e-20, -4.111937e-20, 2.006177e-36, -1.027984e-20, -1.541976e-20, 
    2.006177e-36, 0, 5.139921e-21, -2.055969e-20, 0, -3.597945e-20, 0, 0, 
    1.541976e-20, -1.027984e-20, -2.006177e-36, 1.541976e-20, 1.027984e-20, 
    5.139921e-21, -2.055969e-20, -1.541976e-20, 1.027984e-20, -1.541976e-20, 
    -2.055969e-20, 2.055969e-20, 1.027984e-20, 0, 3.597945e-20, 
    -1.541976e-20, 0, 3.083953e-20, -2.055969e-20, 1.027984e-20, 
    5.139921e-21, 0, 2.006177e-36, -1.541976e-20, 2.055969e-20, 2.055969e-20, 
    -5.139921e-21, -4.625929e-20, 1.541976e-20, 1.541976e-20, -2.055969e-20, 
    -2.569961e-20, 4.111937e-20, 1.027984e-20, 1.541976e-20, 1.541976e-20, 
    1.027984e-20, -5.139921e-21, -1.541976e-20, -4.111937e-20, 5.139921e-21, 
    -5.139921e-21, 0, -5.139921e-21, -1.027984e-20, -5.139921e-21, 
    3.083953e-20, -1.541976e-20, 2.055969e-20, -4.111937e-20, -1.541976e-20, 
    -1.541976e-20, 1.541976e-20, 0, -1.027984e-20, -1.027984e-20, 
    3.597945e-20, 0, -2.055969e-20, -1.541976e-20, 1.027984e-20, 
    -2.055969e-20, 2.569961e-20, 2.006177e-36, 2.569961e-20, 5.139921e-21, 
    1.027984e-20, 0, 1.027984e-20, 3.083953e-20, 2.055969e-20, -2.055969e-20, 
    -3.597945e-20, 2.569961e-20, 0, 1.541976e-20, 2.055969e-20, 
    -1.541976e-20, -5.139921e-21, 5.139921e-21, 0, -5.139921e-21, 0, 
    -5.139921e-21, -1.027984e-20, 1.027984e-20, 5.139921e-21, -1.027984e-20, 
    -2.006177e-36, -5.139921e-21, -1.541976e-20, -1.027984e-20, 5.139921e-21, 
    0, -5.139921e-21, 0, -1.027984e-20, -5.139921e-21, -3.597945e-20, 0, 
    -2.055969e-20, -2.006177e-36, -2.055969e-20, 5.139921e-21, 2.569961e-20, 
    -1.027984e-20, 2.055969e-20, 0, -1.027984e-20, 0, -1.027984e-20, 
    5.139921e-21, 1.541976e-20, -2.006177e-36, -1.027984e-20, 5.139921e-21, 
    5.139921e-21, -1.541976e-20, -2.569961e-20,
  -5.139921e-21, -5.139921e-21, -2.569961e-20, -1.027984e-20, 3.083953e-20, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, -1.027984e-20, -1.541976e-20, 
    -5.139921e-21, 2.569961e-20, 5.139921e-21, 1.027984e-20, -3.083953e-20, 
    -1.027984e-20, -5.139921e-21, 4.111937e-20, -3.083953e-20, 0, 
    -2.006177e-36, 2.055969e-20, 3.083953e-20, 1.027984e-20, -1.541976e-20, 
    -3.597945e-20, -1.541976e-20, 5.139921e-21, 5.139921e-21, -1.541976e-20, 
    5.139921e-21, 1.541976e-20, -5.139921e-21, 1.027984e-20, -1.541976e-20, 
    -1.027984e-20, -1.027984e-20, 0, 0, -5.139921e-21, 0, 5.139921e-21, 
    -5.139921e-21, 0, 5.139921e-21, 1.027984e-20, -1.027984e-20, 0, 0, 
    2.006177e-36, 0, -1.027984e-20, 2.569961e-20, 1.541976e-20, 0, 
    1.541976e-20, 2.055969e-20, -2.569961e-20, -4.111937e-20, 2.055969e-20, 
    1.027984e-20, -3.083953e-20, -5.139921e-21, 0, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 1.541976e-20, -1.027984e-20, -2.006177e-36, 
    -5.139921e-21, -5.139921e-21, 0, 0, -1.541976e-20, 0, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, -1.027984e-20, -1.027984e-20, 2.006177e-36, 
    2.055969e-20, -1.541976e-20, 2.055969e-20, 2.006177e-36, -1.541976e-20, 
    -5.139921e-21, 2.569961e-20, 5.139921e-21, -1.027984e-20, -1.541976e-20, 
    -1.541976e-20, -5.139921e-21, -1.027984e-20, -5.139921e-21, 
    -5.139921e-21, 1.541976e-20, -1.027984e-20, 1.027984e-20, 1.541976e-20, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    -2.055969e-20, 1.027984e-20, 5.139921e-21, 1.541976e-20, -1.541976e-20, 
    -5.139921e-21, 0, 5.139921e-21, -2.569961e-20, 3.597945e-20, 
    -2.055969e-20, -5.139921e-21, -5.139921e-21, 0, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, 0, -1.541976e-20, -5.139921e-21, 
    -1.541976e-20, 1.027984e-20, -1.541976e-20, 5.139921e-21, -5.139921e-21, 
    -1.027984e-20, -1.027984e-20, 1.027984e-20, -1.541976e-20, 1.541976e-20, 
    2.055969e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    0, 2.055969e-20, 2.055969e-20, 1.541976e-20, 5.139921e-21, 5.139921e-21, 
    0, 1.027984e-20, 3.083953e-20, 5.139921e-21, 1.541976e-20, 3.597945e-20, 
    -5.139921e-21, 0, -5.139921e-21, -1.027984e-20, 3.083953e-20, 0, 
    1.027984e-20, -2.006177e-36, -1.541976e-20, 5.139921e-21, 5.139921e-21, 
    5.139921e-21, 1.541976e-20, 2.055969e-20, 0, -1.027984e-20, 
    -1.541976e-20, 5.139921e-21, -5.139921e-21, 0, -1.541976e-20, 
    -5.139921e-21, 5.139921e-21, 1.027984e-20, 0, 3.083953e-20, 0, 
    -5.139921e-21, -2.569961e-20, 2.006177e-36, -2.055969e-20, 1.541976e-20, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, -1.027984e-20, -3.083953e-20, 
    2.006177e-36, -1.027984e-20, 2.055969e-20, -2.055969e-20, -2.055969e-20, 
    5.139921e-21, 5.139921e-21, -5.139921e-21, 1.541976e-20, 1.027984e-20, 
    5.139921e-21, -1.541976e-20, -2.055969e-20, -2.569961e-20, 1.541976e-20, 
    5.139921e-21, 1.541976e-20, 2.055969e-20, -1.541976e-20, -1.541976e-20, 
    -1.027984e-20, -2.006177e-36, 2.569961e-20, -5.139921e-21, -1.027984e-20, 
    1.027984e-20, -1.027984e-20, -5.139921e-21, 5.139921e-21, 1.027984e-20, 
    1.541976e-20, -1.541976e-20, -5.139921e-21, 1.027984e-20, -1.027984e-20, 
    0, -1.027984e-20, 2.006177e-36, 1.027984e-20, 5.139921e-21, 
    -2.055969e-20, 0, 1.541976e-20, -1.541976e-20, 0, 2.006177e-36, 
    1.541976e-20, 5.139921e-21, -5.139921e-21, 0, 1.027984e-20, 
    -1.541976e-20, -1.027984e-20, -2.055969e-20, -3.083953e-20, 
    -5.139921e-21, -3.597945e-20, -1.541976e-20, -2.055969e-20, 1.027984e-20, 
    -1.541976e-20, 1.027984e-20, -5.139921e-21, -5.139921e-21, 1.541976e-20, 
    1.027984e-20, 2.006177e-36, -2.055969e-20, 2.055969e-20, 1.027984e-20, 
    -2.055969e-20, 0, 2.569961e-20, 1.027984e-20, 1.541976e-20, 
    -2.055969e-20, -2.006177e-36, 5.139921e-21, -2.055969e-20, 1.027984e-20, 
    -2.569961e-20, -2.569961e-20, -1.541976e-20, -1.027984e-20, 
    -1.027984e-20, 0, 1.027984e-20, 0, -1.541976e-20, 2.569961e-20, 
    1.541976e-20, 1.027984e-20, -5.139921e-21, -3.083953e-20, 1.027984e-20, 
    0, 1.027984e-20, 5.139921e-21, 1.027984e-20, 5.139921e-21, -1.541976e-20, 
    1.027984e-20, -1.027984e-20, 2.569961e-20, 5.139921e-21, 0, 2.006177e-36, 
    1.541976e-20, 1.541976e-20, 1.027984e-20, 0, -1.541976e-20, 0, 
    -2.055969e-20, 3.083953e-20, -1.541976e-20, 1.027984e-20, 0, 
    -5.139921e-21, 1.027984e-20, 3.083953e-20, -1.541976e-20, 0, 
    2.055969e-20, 1.541976e-20, -2.569961e-20, 5.139921e-21, -1.027984e-20, 
    -1.027984e-20, -1.541976e-20, 5.139921e-21, -2.055969e-20, 2.006177e-36, 
    -1.541976e-20, 1.541976e-20, 1.541976e-20, 1.027984e-20, 1.541976e-20, 
    1.541976e-20, -5.139921e-21, -1.541976e-20, 0, 2.006177e-36, 
    2.055969e-20, 5.139921e-21, 1.027984e-20, -3.597945e-20, -5.139921e-21,
  2.055969e-20, 2.055969e-20, -5.139921e-21, 4.111937e-20, -2.055969e-20, 
    5.139921e-21, -3.083953e-20, -2.569961e-20, -5.139921e-21, -2.569961e-20, 
    1.541976e-20, 5.139921e-21, 1.541976e-20, -5.139921e-21, -1.027984e-20, 
    -1.027984e-20, 5.139921e-21, 1.541976e-20, 1.027984e-20, 0, 
    -2.006177e-36, -1.541976e-20, -1.541976e-20, 0, 0, -1.027984e-20, 
    1.027984e-20, 1.027984e-20, -5.139921e-21, 1.027984e-20, -2.055969e-20, 
    2.055969e-20, 5.139921e-21, -5.139921e-21, 0, -2.055969e-20, 
    -1.027984e-20, -1.027984e-20, 1.027984e-20, -1.027984e-20, 5.139921e-21, 
    -2.055969e-20, 1.027984e-20, 2.569961e-20, 1.027984e-20, -3.597945e-20, 
    0, 0, -1.541976e-20, 2.006177e-36, 5.139921e-21, -5.139921e-21, 
    1.027984e-20, -1.027984e-20, -1.541976e-20, 1.541976e-20, -5.139921e-21, 
    5.139921e-21, 5.139921e-21, -1.541976e-20, 5.139921e-21, -1.541976e-20, 
    -2.055969e-20, 7.19589e-20, 2.569961e-20, 0, 5.139921e-21, 1.027984e-20, 
    -1.027984e-20, -2.055969e-20, -3.083953e-20, -1.027984e-20, 
    -2.055969e-20, 2.569961e-20, 1.541976e-20, 2.055969e-20, 2.569961e-20, 
    1.027984e-20, 0, 5.139921e-21, 5.139921e-20, 3.083953e-20, 5.139921e-21, 
    2.006177e-36, -1.541976e-20, -1.027984e-20, 2.569961e-20, -1.541976e-20, 
    -3.597945e-20, -3.083953e-20, -1.541976e-20, -2.569961e-20, 
    -5.139921e-21, -1.541976e-20, -2.055969e-20, 5.139921e-21, 5.139921e-21, 
    5.139921e-21, 0, -1.027984e-20, 3.083953e-20, 5.139921e-21, 
    -4.625929e-20, 0, -1.027984e-20, 2.055969e-20, 0, -1.541976e-20, 
    2.055969e-20, 5.139921e-21, 2.569961e-20, -5.139921e-21, 2.055969e-20, 
    2.569961e-20, -1.541976e-20, -5.139921e-21, -4.111937e-20, 0, 0, 
    2.055969e-20, -3.083953e-20, 0, -2.006177e-36, 5.139921e-21, 
    -5.139921e-21, 1.027984e-20, 2.569961e-20, 4.111937e-20, 5.139921e-21, 
    -2.569961e-20, 0, -3.083953e-20, -2.055969e-20, -5.139921e-21, 
    1.027984e-20, 0, 2.055969e-20, -1.027984e-20, 2.055969e-20, 
    -2.055969e-20, 2.569961e-20, -5.139921e-21, -1.541976e-20, 1.027984e-20, 
    -2.055969e-20, -5.139921e-21, -2.055969e-20, -2.006177e-36, 2.055969e-20, 
    -1.541976e-20, 2.055969e-20, 5.139921e-21, -2.055969e-20, -1.027984e-20, 
    -2.055969e-20, -1.027984e-20, -1.541976e-20, 1.027984e-20, 2.006177e-36, 
    -2.055969e-20, 5.139921e-21, 1.027984e-20, 5.139921e-21, 3.083953e-20, 
    -1.027984e-20, -1.027984e-20, 1.027984e-20, 1.541976e-20, 5.139921e-21, 
    5.139921e-21, 0, -1.541976e-20, 5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 3.083953e-20, 5.139921e-21, -2.055969e-20, 1.027984e-20, 
    5.139921e-21, -1.541976e-20, 2.569961e-20, -5.139921e-21, 3.083953e-20, 
    2.055969e-20, 3.083953e-20, 1.541976e-20, 2.569961e-20, 1.541976e-20, 
    -1.027984e-20, 0, -1.541976e-20, -5.139921e-21, -5.139921e-21, 
    1.541976e-20, -1.541976e-20, 1.541976e-20, 1.541976e-20, -1.541976e-20, 
    1.027984e-20, 5.139921e-21, 2.055969e-20, -3.597945e-20, 1.541976e-20, 
    -1.027984e-20, -1.027984e-20, 5.139921e-21, -5.139921e-21, 4.111937e-20, 
    -1.027984e-20, 2.006177e-36, 1.541976e-20, 5.139921e-21, 5.139921e-21, 
    2.569961e-20, -5.139921e-21, 3.083953e-20, 1.027984e-20, 2.055969e-20, 
    1.541976e-20, -3.083953e-20, -5.139921e-21, -3.597945e-20, 1.541976e-20, 
    -5.139921e-21, 2.055969e-20, -5.139921e-21, -1.027984e-20, -5.139921e-21, 
    5.139921e-21, -1.027984e-20, -1.541976e-20, 0, -5.139921e-21, 
    -5.139921e-21, 5.139921e-21, -1.027984e-20, -5.139921e-21, 5.139921e-21, 
    -3.083953e-20, 2.055969e-20, -5.139921e-21, -1.027984e-20, -1.541976e-20, 
    -1.541976e-20, 5.139921e-21, -5.139921e-21, -2.055969e-20, 5.139921e-21, 
    -5.139921e-21, 1.541976e-20, -1.541976e-20, -1.027984e-20, 3.083953e-20, 
    -2.055969e-20, 1.027984e-20, -2.055969e-20, 1.541976e-20, -2.569961e-20, 
    -5.139921e-21, 3.597945e-20, 1.541976e-20, -1.027984e-20, -3.083953e-20, 
    5.139921e-21, 3.083953e-20, 2.569961e-20, 1.541976e-20, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, -1.541976e-20, 2.055969e-20, 2.055969e-20, 
    2.569961e-20, -1.541976e-20, 2.569961e-20, 3.597945e-20, 3.083953e-20, 
    1.541976e-20, 1.541976e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    2.055969e-20, -4.111937e-20, 2.006177e-36, 0, -2.569961e-20, 
    1.027984e-20, 5.139921e-21, 5.139921e-21, 0, -1.027984e-20, 1.541976e-20, 
    1.027984e-20, -2.006177e-36, 2.055969e-20, -4.625929e-20, -1.027984e-20, 
    0, -1.027984e-20, -5.139921e-21, -1.027984e-20, -5.139921e-21, 
    -2.006177e-36, 0, 5.139921e-21, -1.541976e-20, -1.027984e-20, 
    2.055969e-20, 1.027984e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    2.055969e-20, -1.541976e-20, 1.541976e-20, 3.083953e-20, -3.083953e-20, 
    -5.139921e-21, -1.027984e-20, 2.006177e-36, -2.055969e-20, 1.027984e-20, 
    -5.139921e-21, 2.055969e-20, -2.055969e-20, 0, -5.139921e-21, 
    -1.541976e-20, 0, 3.083953e-20, -5.139921e-21, 2.569961e-20, 0, 
    1.027984e-20, 2.055969e-20,
  2.055969e-20, -5.139921e-21, 5.139921e-21, 1.541976e-20, 5.139921e-21, 
    -5.139921e-21, 2.055969e-20, 5.139921e-21, 0, 0, -2.055969e-20, 
    -5.139921e-21, -1.541976e-20, 3.083953e-20, -1.541976e-20, 1.027984e-20, 
    2.055969e-20, -1.027984e-20, -1.541976e-20, 2.055969e-20, -3.597945e-20, 
    1.027984e-20, 0, -2.569961e-20, -5.139921e-21, -5.139921e-21, 
    -1.541976e-20, 1.027984e-20, -1.541976e-20, -1.541976e-20, 1.027984e-20, 
    -1.541976e-20, 3.083953e-20, 1.541976e-20, -1.027984e-20, 2.006177e-36, 
    1.027984e-20, -5.139921e-21, -1.027984e-20, 2.569961e-20, -1.541976e-20, 
    2.055969e-20, -2.006177e-36, 2.055969e-20, 1.027984e-20, 1.541976e-20, 
    -1.027984e-20, 4.111937e-20, 1.541976e-20, 2.569961e-20, -5.139921e-21, 
    -3.083953e-20, 0, -3.083953e-20, -1.541976e-20, 5.139921e-21, 
    -5.139921e-21, -2.569961e-20, -3.083953e-20, 1.027984e-20, 0, 
    3.597945e-20, -5.139921e-21, -3.083953e-20, -2.055969e-20, -1.541976e-20, 
    -1.027984e-20, 5.139921e-21, -5.139921e-21, -2.055969e-20, 1.027984e-20, 
    -1.541976e-20, -2.055969e-20, 2.055969e-20, -5.139921e-21, -1.027984e-20, 
    -1.027984e-20, -2.006177e-36, -2.006177e-36, -5.139921e-21, 1.541976e-20, 
    1.541976e-20, 1.541976e-20, 1.027984e-20, -2.055969e-20, 2.569961e-20, 
    1.027984e-20, -2.055969e-20, 1.541976e-20, -1.541976e-20, -4.111937e-20, 
    2.055969e-20, -2.055969e-20, 2.569961e-20, 5.139921e-21, 5.139921e-21, 
    1.027984e-20, -2.055969e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -5.139921e-20, 1.027984e-20, 1.027984e-20, 1.541976e-20, -2.055969e-20, 
    1.027984e-20, 5.139921e-21, 1.027984e-20, 0, -3.083953e-20, 4.111937e-20, 
    1.027984e-20, -1.027984e-20, -5.139921e-21, -3.083953e-20, -2.569961e-20, 
    2.569961e-20, 3.083953e-20, 1.541976e-20, 2.055969e-20, 5.139921e-21, 
    5.139921e-21, 2.569961e-20, 2.006177e-36, 5.139921e-21, 0, 0, 
    1.541976e-20, 1.027984e-20, -1.541976e-20, 2.569961e-20, -1.541976e-20, 
    -3.083953e-20, 5.139921e-21, 1.027984e-20, -1.027984e-20, -5.139921e-21, 
    1.541976e-20, -1.541976e-20, -1.027984e-20, -3.597945e-20, -3.083953e-20, 
    -4.111937e-20, 5.139921e-21, 2.006177e-36, 2.569961e-20, -1.541976e-20, 
    2.055969e-20, 3.083953e-20, -3.083953e-20, -1.541976e-20, -5.139921e-21, 
    2.006177e-36, -2.006177e-36, 1.541976e-20, -3.597945e-20, 2.055969e-20, 
    3.083953e-20, -2.006177e-36, 0, -2.055969e-20, -3.083953e-20, 
    2.006177e-36, 0, 5.139921e-20, -5.139921e-21, 3.597945e-20, 1.541976e-20, 
    -3.083953e-20, 3.597945e-20, -2.055969e-20, 5.139921e-21, 0, 
    -5.139921e-21, -1.541976e-20, -1.541976e-20, -5.139921e-21, 4.625929e-20, 
    -3.083953e-20, 0, -2.055969e-20, -1.541976e-20, 0, -1.027984e-20, 
    -2.055969e-20, -5.139921e-21, -3.597945e-20, -3.083953e-20, 1.541976e-20, 
    2.006177e-36, 5.139921e-21, 2.055969e-20, 2.055969e-20, -3.597945e-20, 
    -5.139921e-21, 5.139921e-21, 0, -5.139921e-21, -2.006177e-36, 0, 
    -2.569961e-20, 3.083953e-20, 3.597945e-20, 0, 2.569961e-20, 2.569961e-20, 
    3.597945e-20, -1.027984e-20, 2.006177e-36, -2.055969e-20, 5.139921e-21, 
    2.569961e-20, -1.541976e-20, 2.006177e-36, 0, 5.139921e-21, 
    -4.111937e-20, -1.541976e-20, -3.083953e-20, -1.027984e-20, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 0, -5.139921e-21, -2.055969e-20, 
    5.139921e-21, -4.111937e-20, -3.083953e-20, -1.541976e-20, -2.569961e-20, 
    2.006177e-36, 5.139921e-21, -1.541976e-20, -1.541976e-20, -4.625929e-20, 
    -5.139921e-21, -5.139921e-21, -1.541976e-20, 0, -1.541976e-20, 
    5.139921e-21, 2.055969e-20, -5.139921e-21, -5.139921e-21, 0, 0, 
    -3.597945e-20, 2.055969e-20, -2.055969e-20, -2.569961e-20, 0, 
    5.139921e-21, -1.027984e-20, 2.006177e-36, -2.055969e-20, -1.027984e-20, 
    -5.139921e-21, -2.055969e-20, 5.139921e-21, 2.569961e-20, -1.027984e-20, 
    1.541976e-20, -1.541976e-20, 1.027984e-20, -4.625929e-20, 5.139921e-21, 
    -4.625929e-20, 2.569961e-20, 4.111937e-20, 5.139921e-21, -1.027984e-20, 
    -2.055969e-20, -1.027984e-20, -1.541976e-20, -2.055969e-20, 
    -3.083953e-20, -3.597945e-20, -1.027984e-20, 3.083953e-20, 2.055969e-20, 
    3.083953e-20, -5.139921e-21, -2.569961e-20, 1.541976e-20, -2.055969e-20, 
    -2.055969e-20, 3.083953e-20, 2.569961e-20, 3.083953e-20, -5.139921e-21, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, -5.139921e-21, 1.541976e-20, 
    -1.541976e-20, -1.541976e-20, 0, -2.055969e-20, 0, -5.139921e-21, 0, 
    5.139921e-21, -1.027984e-20, 2.569961e-20, -2.569961e-20, -3.597945e-20, 
    -2.055969e-20, -5.139921e-21, 4.625929e-20, 1.027984e-20, 3.597945e-20, 
    -1.541976e-20, 1.027984e-20, -2.006177e-36, -1.027984e-20, 5.139921e-21, 
    2.055969e-20, 1.541976e-20, -1.541976e-20, 5.139921e-21, -1.541976e-20, 
    -5.139921e-21, -5.139921e-21, 2.569961e-20, -2.055969e-20, 3.597945e-20, 
    5.139921e-21, -2.006177e-36, 5.139921e-21, 5.139921e-21, -1.027984e-20, 
    2.006177e-36, 5.139921e-20, 5.139921e-21, -1.027984e-20,
  3.083953e-20, -1.541976e-20, -1.027984e-20, -1.027984e-20, -2.006177e-36, 
    -2.569961e-20, 2.569961e-20, 1.027984e-20, -1.541976e-20, -5.139921e-21, 
    0, 0, 1.541976e-20, -1.027984e-20, 5.139921e-21, 2.006177e-36, 0, 0, 
    -2.055969e-20, 0, 5.139921e-21, 5.139921e-21, 0, 0, -5.139921e-21, 
    1.027984e-20, 2.006177e-36, -5.139921e-21, 3.083953e-20, -1.027984e-20, 
    -5.139921e-21, -3.597945e-20, -2.569961e-20, 1.027984e-20, 1.541976e-20, 
    1.541976e-20, 1.541976e-20, 1.027984e-20, -2.055969e-20, 2.055969e-20, 0, 
    1.027984e-20, 5.139921e-21, 2.569961e-20, 1.027984e-20, 1.027984e-20, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, 5.139921e-21, -1.541976e-20, 
    2.055969e-20, 0, 1.027984e-20, 2.055969e-20, 1.541976e-20, -5.139921e-21, 
    1.541976e-20, 1.541976e-20, 5.139921e-21, -2.055969e-20, 2.055969e-20, 
    5.139921e-21, 5.139921e-21, -1.027984e-20, 3.083953e-20, -1.027984e-20, 
    1.541976e-20, 4.625929e-20, -2.055969e-20, 3.083953e-20, 1.027984e-20, 
    2.006177e-36, 5.139921e-21, -1.541976e-20, -1.027984e-20, 2.569961e-20, 
    2.055969e-20, 1.027984e-20, -1.541976e-20, 1.541976e-20, -3.083953e-20, 
    -4.625929e-20, 1.541976e-20, -2.569961e-20, -2.055969e-20, 1.541976e-20, 
    0, 2.569961e-20, -3.083953e-20, 0, 5.139921e-21, 1.541976e-20, 
    -2.569961e-20, -2.055969e-20, 1.027984e-20, -3.083953e-20, 1.027984e-20, 
    -5.139921e-21, 1.541976e-20, -1.027984e-20, -2.055969e-20, 5.139921e-21, 
    -5.139921e-21, -1.027984e-20, -4.625929e-20, 1.027984e-20, 1.027984e-20, 
    1.541976e-20, -1.541976e-20, 2.569961e-20, -1.027984e-20, -1.541976e-20, 
    -1.541976e-20, 1.541976e-20, 3.597945e-20, 0, 5.139921e-21, 1.027984e-20, 
    1.027984e-20, -2.569961e-20, 2.569961e-20, 5.139921e-21, 1.027984e-20, 
    2.006177e-36, 2.569961e-20, 1.541976e-20, 2.055969e-20, 1.541976e-20, 
    -1.541976e-20, 5.139921e-21, 5.139921e-21, -3.597945e-20, -5.139921e-21, 
    -2.569961e-20, 0, -3.597945e-20, -3.083953e-20, 5.139921e-21, 
    3.083953e-20, 0, 5.139921e-21, 3.083953e-20, 0, 2.055969e-20, 
    5.139921e-21, -1.541976e-20, 2.055969e-20, -3.083953e-20, 0, 
    -2.006177e-36, -2.569961e-20, -1.027984e-20, -5.139921e-21, 
    -1.027984e-20, 2.055969e-20, -1.027984e-20, 2.055969e-20, 5.139921e-21, 
    -3.597945e-20, -5.139921e-21, -5.139921e-21, 3.597945e-20, -1.541976e-20, 
    1.027984e-20, -4.625929e-20, 5.139921e-21, -5.139921e-20, 2.006177e-36, 
    5.139921e-21, 5.139921e-21, 1.027984e-20, 2.569961e-20, 1.027984e-20, 
    -2.055969e-20, 3.083953e-20, 2.055969e-20, -2.006177e-36, 1.027984e-20, 
    1.027984e-20, -2.569961e-20, 5.139921e-21, -1.541976e-20, -1.027984e-20, 
    -2.055969e-20, 5.139921e-21, -2.006177e-36, 2.569961e-20, 5.139921e-21, 
    -2.569961e-20, 4.111937e-20, -1.541976e-20, 2.055969e-20, -1.541976e-20, 
    0, 2.569961e-20, -5.139921e-21, 1.027984e-20, 2.055969e-20, 
    -1.027984e-20, 2.569961e-20, 1.027984e-20, 1.027984e-20, 1.027984e-20, 
    3.597945e-20, -2.569961e-20, 2.055969e-20, 5.139921e-21, -2.569961e-20, 
    -5.139921e-21, 1.541976e-20, -2.006177e-36, -1.541976e-20, 2.006177e-36, 
    -2.055969e-20, 2.006177e-36, -1.027984e-20, 2.055969e-20, 2.569961e-20, 
    3.083953e-20, 1.027984e-20, -5.139921e-21, 0, 1.541976e-20, 1.027984e-20, 
    -5.139921e-21, -1.541976e-20, -2.569961e-20, 0, 5.139921e-21, 
    5.139921e-21, -2.055969e-20, 1.027984e-20, -1.027984e-20, 1.027984e-20, 
    1.541976e-20, -2.055969e-20, 0, -2.006177e-36, 1.541976e-20, 
    -2.569961e-20, 1.541976e-20, 3.083953e-20, 5.139921e-21, -2.055969e-20, 
    -1.541976e-20, -1.027984e-20, 5.139921e-21, -1.541976e-20, 1.541976e-20, 
    2.055969e-20, 1.541976e-20, -4.111937e-20, -1.541976e-20, -5.139921e-21, 
    4.111937e-20, 5.139921e-21, -1.027984e-20, -3.083953e-20, -1.027984e-20, 
    -5.139921e-21, -3.597945e-20, -1.541976e-20, 5.139921e-21, -1.027984e-20, 
    -2.569961e-20, 1.027984e-20, -1.027984e-20, 5.139921e-21, -1.027984e-20, 
    -1.027984e-20, 0, 5.139921e-21, 1.027984e-20, 3.083953e-20, 
    -2.569961e-20, -1.541976e-20, 1.027984e-20, 1.541976e-20, 5.139921e-21, 
    0, -1.027984e-20, 4.625929e-20, 1.027984e-20, -1.541976e-20, 
    -2.055969e-20, 2.569961e-20, -1.027984e-20, 1.541976e-20, 5.139921e-21, 
    2.569961e-20, 1.541976e-20, 3.597945e-20, -1.027984e-20, -1.027984e-20, 
    -2.055969e-20, -2.006177e-36, -1.027984e-20, 0, 2.006177e-36, 
    -1.541976e-20, 0, -1.027984e-20, 1.027984e-20, 2.569961e-20, 
    2.055969e-20, -5.139921e-21, 1.541976e-20, -5.139921e-21, 2.055969e-20, 
    1.541976e-20, -1.027984e-20, -1.541976e-20, 1.027984e-20, -2.055969e-20, 
    5.139921e-21, -1.541976e-20, -1.541976e-20, 1.027984e-20, 3.083953e-20, 
    -3.597945e-20, 5.139921e-21, -1.027984e-20, -2.055969e-20, 2.055969e-20, 
    1.027984e-20, 1.541976e-20, -5.139921e-21, -5.139921e-21, 1.541976e-20, 
    0, 2.006177e-36, 3.597945e-20, -1.541976e-20, -1.541976e-20, 
    2.006177e-36, 1.541976e-20, 2.055969e-20,
  8.598664e-29, 8.598635e-29, 8.598641e-29, 8.598618e-29, 8.59863e-29, 
    8.598615e-29, 8.598658e-29, 8.598634e-29, 8.598649e-29, 8.598662e-29, 
    8.598573e-29, 8.598617e-29, 8.598527e-29, 8.598556e-29, 8.598485e-29, 
    8.598532e-29, 8.598476e-29, 8.598486e-29, 8.598454e-29, 8.598463e-29, 
    8.598422e-29, 8.59845e-29, 8.5984e-29, 8.598429e-29, 8.598424e-29, 
    8.598451e-29, 8.598608e-29, 8.598578e-29, 8.59861e-29, 8.598606e-29, 
    8.598607e-29, 8.59863e-29, 8.598642e-29, 8.598666e-29, 8.598662e-29, 
    8.598644e-29, 8.598604e-29, 8.598617e-29, 8.598583e-29, 8.598583e-29, 
    8.598545e-29, 8.598562e-29, 8.598498e-29, 8.598516e-29, 8.598463e-29, 
    8.598476e-29, 8.598463e-29, 8.598468e-29, 8.598463e-29, 8.598483e-29, 
    8.598475e-29, 8.598492e-29, 8.598559e-29, 8.598539e-29, 8.598598e-29, 
    8.598633e-29, 8.598657e-29, 8.598674e-29, 8.598671e-29, 8.598667e-29, 
    8.598643e-29, 8.598622e-29, 8.598606e-29, 8.598595e-29, 8.598584e-29, 
    8.598551e-29, 8.598533e-29, 8.598494e-29, 8.598501e-29, 8.598489e-29, 
    8.598478e-29, 8.598459e-29, 8.598462e-29, 8.598453e-29, 8.598489e-29, 
    8.598465e-29, 8.598505e-29, 8.598494e-29, 8.598581e-29, 8.598613e-29, 
    8.598627e-29, 8.59864e-29, 8.598669e-29, 8.598649e-29, 8.598657e-29, 
    8.598638e-29, 8.598625e-29, 8.598631e-29, 8.598594e-29, 8.598609e-29, 
    8.598532e-29, 8.598565e-29, 8.598479e-29, 8.5985e-29, 8.598474e-29, 
    8.598487e-29, 8.598465e-29, 8.598485e-29, 8.59845e-29, 8.598442e-29, 
    8.598448e-29, 8.598427e-29, 8.598486e-29, 8.598463e-29, 8.598632e-29, 
    8.598631e-29, 8.598626e-29, 8.598646e-29, 8.598648e-29, 8.598666e-29, 
    8.598649e-29, 8.598643e-29, 8.598625e-29, 8.598614e-29, 8.598604e-29, 
    8.598582e-29, 8.598557e-29, 8.598523e-29, 8.598498e-29, 8.598482e-29, 
    8.598492e-29, 8.598483e-29, 8.598493e-29, 8.598498e-29, 8.598445e-29, 
    8.598475e-29, 8.59843e-29, 8.598433e-29, 8.598453e-29, 8.598433e-29, 
    8.59863e-29, 8.598636e-29, 8.598655e-29, 8.59864e-29, 8.598668e-29, 
    8.598652e-29, 8.598643e-29, 8.598609e-29, 8.598601e-29, 8.598593e-29, 
    8.59858e-29, 8.598562e-29, 8.59853e-29, 8.598502e-29, 8.598477e-29, 
    8.598479e-29, 8.598478e-29, 8.598473e-29, 8.598486e-29, 8.59847e-29, 
    8.598468e-29, 8.598475e-29, 8.598433e-29, 8.598445e-29, 8.598433e-29, 
    8.598441e-29, 8.598634e-29, 8.598624e-29, 8.59863e-29, 8.59862e-29, 
    8.598627e-29, 8.598596e-29, 8.598587e-29, 8.598544e-29, 8.598562e-29, 
    8.598534e-29, 8.598559e-29, 8.598554e-29, 8.598533e-29, 8.598557e-29, 
    8.598504e-29, 8.598541e-29, 8.598473e-29, 8.598509e-29, 8.59847e-29, 
    8.598477e-29, 8.598465e-29, 8.598455e-29, 8.598442e-29, 8.598418e-29, 
    8.598423e-29, 8.598403e-29, 8.59861e-29, 8.598598e-29, 8.598599e-29, 
    8.598586e-29, 8.598576e-29, 8.598556e-29, 8.598522e-29, 8.598535e-29, 
    8.598512e-29, 8.598507e-29, 8.598542e-29, 8.59852e-29, 8.598589e-29, 
    8.598578e-29, 8.598585e-29, 8.598609e-29, 8.598532e-29, 8.598571e-29, 
    8.598498e-29, 8.598519e-29, 8.598456e-29, 8.598488e-29, 8.598426e-29, 
    8.5984e-29, 8.598375e-29, 8.598346e-29, 8.598591e-29, 8.5986e-29, 
    8.598584e-29, 8.598563e-29, 8.598544e-29, 8.598518e-29, 8.598515e-29, 
    8.59851e-29, 8.598498e-29, 8.598488e-29, 8.598509e-29, 8.598485e-29, 
    8.598575e-29, 8.598528e-29, 8.598603e-29, 8.59858e-29, 8.598565e-29, 
    8.598571e-29, 8.598536e-29, 8.598527e-29, 8.598494e-29, 8.598511e-29, 
    8.598406e-29, 8.598453e-29, 8.598324e-29, 8.59836e-29, 8.598603e-29, 
    8.598591e-29, 8.598551e-29, 8.59857e-29, 8.598516e-29, 8.598503e-29, 
    8.598492e-29, 8.598479e-29, 8.598477e-29, 8.598469e-29, 8.598482e-29, 
    8.59847e-29, 8.598518e-29, 8.598497e-29, 8.598556e-29, 8.598541e-29, 
    8.598548e-29, 8.598556e-29, 8.598533e-29, 8.598509e-29, 8.598508e-29, 
    8.598501e-29, 8.598479e-29, 8.598516e-29, 8.5984e-29, 8.598472e-29, 
    8.598578e-29, 8.598557e-29, 8.598554e-29, 8.598562e-29, 8.598504e-29, 
    8.598525e-29, 8.598469e-29, 8.598485e-29, 8.598459e-29, 8.598472e-29, 
    8.598474e-29, 8.598489e-29, 8.5985e-29, 8.598524e-29, 8.598545e-29, 
    8.598561e-29, 8.598557e-29, 8.598539e-29, 8.598507e-29, 8.598477e-29, 
    8.598483e-29, 8.598461e-29, 8.59852e-29, 8.598495e-29, 8.598505e-29, 
    8.59848e-29, 8.598535e-29, 8.598488e-29, 8.598547e-29, 8.598542e-29, 
    8.598525e-29, 8.598494e-29, 8.598487e-29, 8.598479e-29, 8.598484e-29, 
    8.598506e-29, 8.59851e-29, 8.598526e-29, 8.59853e-29, 8.598543e-29, 
    8.598553e-29, 8.598544e-29, 8.598534e-29, 8.598506e-29, 8.598482e-29, 
    8.598455e-29, 8.598448e-29, 8.598417e-29, 8.598442e-29, 8.5984e-29, 
    8.598436e-29, 8.598374e-29, 8.598486e-29, 8.598437e-29, 8.598525e-29, 
    8.598516e-29, 8.598498e-29, 8.598459e-29, 8.59848e-29, 8.598456e-29, 
    8.59851e-29, 8.598539e-29, 8.598546e-29, 8.59856e-29, 8.598546e-29, 
    8.598547e-29, 8.598533e-29, 8.598538e-29, 8.598506e-29, 8.598523e-29, 
    8.598474e-29, 8.598456e-29, 8.598405e-29, 8.598374e-29, 8.598342e-29, 
    8.598328e-29, 8.598324e-29, 8.598322e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N_TO_SOIL2N =
  1.164952e-08, 1.170074e-08, 1.169078e-08, 1.173209e-08, 1.170917e-08, 
    1.173622e-08, 1.16599e-08, 1.170277e-08, 1.16754e-08, 1.165413e-08, 
    1.181225e-08, 1.173393e-08, 1.18936e-08, 1.184365e-08, 1.196912e-08, 
    1.188583e-08, 1.198592e-08, 1.196672e-08, 1.20245e-08, 1.200795e-08, 
    1.208186e-08, 1.203214e-08, 1.212017e-08, 1.206998e-08, 1.207783e-08, 
    1.20305e-08, 1.174969e-08, 1.18025e-08, 1.174656e-08, 1.175409e-08, 
    1.175071e-08, 1.170965e-08, 1.168895e-08, 1.16456e-08, 1.165347e-08, 
    1.168531e-08, 1.175748e-08, 1.173298e-08, 1.179472e-08, 1.179333e-08, 
    1.186206e-08, 1.183107e-08, 1.194659e-08, 1.191376e-08, 1.200864e-08, 
    1.198478e-08, 1.200752e-08, 1.200062e-08, 1.200761e-08, 1.197261e-08, 
    1.198761e-08, 1.195681e-08, 1.183687e-08, 1.187212e-08, 1.176699e-08, 
    1.170378e-08, 1.166178e-08, 1.163199e-08, 1.16362e-08, 1.164423e-08, 
    1.16855e-08, 1.172429e-08, 1.175386e-08, 1.177364e-08, 1.179313e-08, 
    1.185211e-08, 1.188333e-08, 1.195323e-08, 1.194062e-08, 1.196199e-08, 
    1.19824e-08, 1.201668e-08, 1.201104e-08, 1.202614e-08, 1.196142e-08, 
    1.200444e-08, 1.193343e-08, 1.195285e-08, 1.179843e-08, 1.173959e-08, 
    1.171458e-08, 1.169269e-08, 1.163944e-08, 1.167621e-08, 1.166172e-08, 
    1.169621e-08, 1.171812e-08, 1.170728e-08, 1.177418e-08, 1.174817e-08, 
    1.188518e-08, 1.182617e-08, 1.198002e-08, 1.194321e-08, 1.198885e-08, 
    1.196556e-08, 1.200546e-08, 1.196955e-08, 1.203176e-08, 1.204531e-08, 
    1.203605e-08, 1.207161e-08, 1.196756e-08, 1.200752e-08, 1.170698e-08, 
    1.170875e-08, 1.171698e-08, 1.168078e-08, 1.167857e-08, 1.164539e-08, 
    1.167491e-08, 1.168748e-08, 1.171939e-08, 1.173827e-08, 1.175621e-08, 
    1.179566e-08, 1.183972e-08, 1.190133e-08, 1.194559e-08, 1.197526e-08, 
    1.195707e-08, 1.197313e-08, 1.195518e-08, 1.194676e-08, 1.204023e-08, 
    1.198775e-08, 1.20665e-08, 1.206214e-08, 1.20265e-08, 1.206263e-08, 
    1.170999e-08, 1.169982e-08, 1.16645e-08, 1.169214e-08, 1.164178e-08, 
    1.166997e-08, 1.168618e-08, 1.174872e-08, 1.176246e-08, 1.17752e-08, 
    1.180036e-08, 1.183266e-08, 1.188931e-08, 1.19386e-08, 1.198359e-08, 
    1.198029e-08, 1.198146e-08, 1.199151e-08, 1.196661e-08, 1.19956e-08, 
    1.200046e-08, 1.198774e-08, 1.206155e-08, 1.204047e-08, 1.206205e-08, 
    1.204831e-08, 1.170312e-08, 1.172024e-08, 1.171099e-08, 1.172838e-08, 
    1.171613e-08, 1.177062e-08, 1.178695e-08, 1.186339e-08, 1.183202e-08, 
    1.188195e-08, 1.183709e-08, 1.184504e-08, 1.188358e-08, 1.183952e-08, 
    1.193588e-08, 1.187055e-08, 1.19919e-08, 1.192666e-08, 1.199599e-08, 
    1.19834e-08, 1.200424e-08, 1.202291e-08, 1.204639e-08, 1.208973e-08, 
    1.207969e-08, 1.211593e-08, 1.174576e-08, 1.176796e-08, 1.176601e-08, 
    1.178924e-08, 1.180642e-08, 1.184366e-08, 1.19034e-08, 1.188093e-08, 
    1.192217e-08, 1.193045e-08, 1.18678e-08, 1.190627e-08, 1.178282e-08, 
    1.180277e-08, 1.179089e-08, 1.174751e-08, 1.188611e-08, 1.181498e-08, 
    1.194633e-08, 1.190779e-08, 1.202025e-08, 1.196432e-08, 1.207417e-08, 
    1.212113e-08, 1.216532e-08, 1.221697e-08, 1.178008e-08, 1.176499e-08, 
    1.1792e-08, 1.182937e-08, 1.186405e-08, 1.191014e-08, 1.191486e-08, 
    1.19235e-08, 1.194586e-08, 1.196467e-08, 1.192623e-08, 1.196939e-08, 
    1.180739e-08, 1.189229e-08, 1.175929e-08, 1.179934e-08, 1.182717e-08, 
    1.181496e-08, 1.187837e-08, 1.189331e-08, 1.195404e-08, 1.192265e-08, 
    1.210954e-08, 1.202685e-08, 1.225629e-08, 1.219217e-08, 1.175972e-08, 
    1.178002e-08, 1.185069e-08, 1.181707e-08, 1.191322e-08, 1.193689e-08, 
    1.195613e-08, 1.198072e-08, 1.198338e-08, 1.199795e-08, 1.197407e-08, 
    1.199701e-08, 1.191024e-08, 1.194902e-08, 1.184261e-08, 1.186851e-08, 
    1.18566e-08, 1.184353e-08, 1.188386e-08, 1.192683e-08, 1.192775e-08, 
    1.194153e-08, 1.198036e-08, 1.191361e-08, 1.212021e-08, 1.199262e-08, 
    1.180217e-08, 1.184128e-08, 1.184686e-08, 1.183171e-08, 1.193452e-08, 
    1.189727e-08, 1.199759e-08, 1.197048e-08, 1.201491e-08, 1.199283e-08, 
    1.198958e-08, 1.196123e-08, 1.194357e-08, 1.189897e-08, 1.186269e-08, 
    1.183391e-08, 1.18406e-08, 1.187221e-08, 1.192946e-08, 1.198362e-08, 
    1.197176e-08, 1.201153e-08, 1.190625e-08, 1.19504e-08, 1.193333e-08, 
    1.197782e-08, 1.188034e-08, 1.196336e-08, 1.185912e-08, 1.186826e-08, 
    1.189653e-08, 1.195339e-08, 1.196597e-08, 1.19794e-08, 1.197111e-08, 
    1.193091e-08, 1.192433e-08, 1.189584e-08, 1.188797e-08, 1.186627e-08, 
    1.18483e-08, 1.186472e-08, 1.188196e-08, 1.193093e-08, 1.197506e-08, 
    1.202317e-08, 1.203495e-08, 1.209117e-08, 1.20454e-08, 1.212092e-08, 
    1.205672e-08, 1.216786e-08, 1.196817e-08, 1.205483e-08, 1.189781e-08, 
    1.191473e-08, 1.194533e-08, 1.20155e-08, 1.197761e-08, 1.202192e-08, 
    1.192407e-08, 1.18733e-08, 1.186016e-08, 1.183566e-08, 1.186072e-08, 
    1.185869e-08, 1.188267e-08, 1.187497e-08, 1.193256e-08, 1.190162e-08, 
    1.19895e-08, 1.202157e-08, 1.211213e-08, 1.216765e-08, 1.222416e-08, 
    1.224911e-08, 1.22567e-08, 1.225988e-08 ;

 SOIL1N_TO_SOIL3N =
  1.382178e-10, 1.388257e-10, 1.387075e-10, 1.391978e-10, 1.389258e-10, 
    1.392469e-10, 1.38341e-10, 1.388498e-10, 1.38525e-10, 1.382725e-10, 
    1.401493e-10, 1.392197e-10, 1.411149e-10, 1.40522e-10, 1.420113e-10, 
    1.410226e-10, 1.422107e-10, 1.419828e-10, 1.426686e-10, 1.424721e-10, 
    1.433494e-10, 1.427593e-10, 1.438042e-10, 1.432085e-10, 1.433017e-10, 
    1.427399e-10, 1.394067e-10, 1.400336e-10, 1.393696e-10, 1.39459e-10, 
    1.394189e-10, 1.389314e-10, 1.386858e-10, 1.381713e-10, 1.382647e-10, 
    1.386426e-10, 1.394992e-10, 1.392084e-10, 1.399412e-10, 1.399247e-10, 
    1.407405e-10, 1.403727e-10, 1.417439e-10, 1.413542e-10, 1.424803e-10, 
    1.421971e-10, 1.424671e-10, 1.423852e-10, 1.424681e-10, 1.420527e-10, 
    1.422307e-10, 1.418652e-10, 1.404415e-10, 1.4086e-10, 1.396121e-10, 
    1.388618e-10, 1.383633e-10, 1.380097e-10, 1.380597e-10, 1.38155e-10, 
    1.386448e-10, 1.391053e-10, 1.394562e-10, 1.39691e-10, 1.399223e-10, 
    1.406224e-10, 1.40993e-10, 1.418227e-10, 1.41673e-10, 1.419266e-10, 
    1.421689e-10, 1.425758e-10, 1.425088e-10, 1.426881e-10, 1.419199e-10, 
    1.424305e-10, 1.415877e-10, 1.418182e-10, 1.399852e-10, 1.392868e-10, 
    1.3899e-10, 1.387302e-10, 1.380981e-10, 1.385346e-10, 1.383626e-10, 
    1.387719e-10, 1.39032e-10, 1.389034e-10, 1.396974e-10, 1.393887e-10, 
    1.410149e-10, 1.403145e-10, 1.421407e-10, 1.417037e-10, 1.422454e-10, 
    1.41969e-10, 1.424427e-10, 1.420164e-10, 1.427548e-10, 1.429156e-10, 
    1.428057e-10, 1.432278e-10, 1.419927e-10, 1.424671e-10, 1.388998e-10, 
    1.389208e-10, 1.390185e-10, 1.385888e-10, 1.385626e-10, 1.381688e-10, 
    1.385192e-10, 1.386684e-10, 1.390471e-10, 1.392712e-10, 1.394841e-10, 
    1.399524e-10, 1.404754e-10, 1.412067e-10, 1.41732e-10, 1.420842e-10, 
    1.418682e-10, 1.420589e-10, 1.418458e-10, 1.417459e-10, 1.428554e-10, 
    1.422324e-10, 1.431671e-10, 1.431154e-10, 1.426924e-10, 1.431212e-10, 
    1.389355e-10, 1.388148e-10, 1.383955e-10, 1.387236e-10, 1.381259e-10, 
    1.384605e-10, 1.386529e-10, 1.393952e-10, 1.395583e-10, 1.397095e-10, 
    1.400082e-10, 1.403915e-10, 1.410639e-10, 1.41649e-10, 1.42183e-10, 
    1.421439e-10, 1.421577e-10, 1.42277e-10, 1.419815e-10, 1.423255e-10, 
    1.423833e-10, 1.422323e-10, 1.431085e-10, 1.428581e-10, 1.431143e-10, 
    1.429513e-10, 1.38854e-10, 1.390572e-10, 1.389474e-10, 1.391538e-10, 
    1.390084e-10, 1.396551e-10, 1.39849e-10, 1.407563e-10, 1.403839e-10, 
    1.409765e-10, 1.404441e-10, 1.405385e-10, 1.409959e-10, 1.404729e-10, 
    1.416167e-10, 1.408413e-10, 1.422816e-10, 1.415073e-10, 1.423302e-10, 
    1.421807e-10, 1.424281e-10, 1.426497e-10, 1.429285e-10, 1.434429e-10, 
    1.433238e-10, 1.437539e-10, 1.393601e-10, 1.396236e-10, 1.396004e-10, 
    1.398762e-10, 1.400801e-10, 1.405221e-10, 1.412311e-10, 1.409645e-10, 
    1.41454e-10, 1.415522e-10, 1.408086e-10, 1.412652e-10, 1.397999e-10, 
    1.400367e-10, 1.398957e-10, 1.393809e-10, 1.41026e-10, 1.401817e-10, 
    1.417407e-10, 1.412833e-10, 1.426181e-10, 1.419543e-10, 1.432582e-10, 
    1.438156e-10, 1.443402e-10, 1.449533e-10, 1.397674e-10, 1.395883e-10, 
    1.399089e-10, 1.403525e-10, 1.407641e-10, 1.413112e-10, 1.413672e-10, 
    1.414697e-10, 1.417352e-10, 1.419584e-10, 1.415021e-10, 1.420144e-10, 
    1.400916e-10, 1.410993e-10, 1.395207e-10, 1.39996e-10, 1.403264e-10, 
    1.401814e-10, 1.409341e-10, 1.411114e-10, 1.418323e-10, 1.414596e-10, 
    1.43678e-10, 1.426965e-10, 1.4542e-10, 1.446589e-10, 1.395258e-10, 
    1.397668e-10, 1.406056e-10, 1.402065e-10, 1.413478e-10, 1.416287e-10, 
    1.41857e-10, 1.42149e-10, 1.421805e-10, 1.423535e-10, 1.4207e-10, 
    1.423423e-10, 1.413124e-10, 1.417726e-10, 1.405097e-10, 1.408171e-10, 
    1.406757e-10, 1.405205e-10, 1.409993e-10, 1.415093e-10, 1.415202e-10, 
    1.416837e-10, 1.421447e-10, 1.413524e-10, 1.438048e-10, 1.422903e-10, 
    1.400296e-10, 1.404938e-10, 1.405601e-10, 1.403803e-10, 1.416005e-10, 
    1.411584e-10, 1.423492e-10, 1.420274e-10, 1.425547e-10, 1.422927e-10, 
    1.422541e-10, 1.419176e-10, 1.41708e-10, 1.411787e-10, 1.407479e-10, 
    1.404063e-10, 1.404858e-10, 1.40861e-10, 1.415405e-10, 1.421834e-10, 
    1.420425e-10, 1.425147e-10, 1.41265e-10, 1.41789e-10, 1.415865e-10, 
    1.421146e-10, 1.409574e-10, 1.419429e-10, 1.407056e-10, 1.408141e-10, 
    1.411496e-10, 1.418246e-10, 1.419739e-10, 1.421333e-10, 1.420349e-10, 
    1.415578e-10, 1.414796e-10, 1.411414e-10, 1.410481e-10, 1.407904e-10, 
    1.405771e-10, 1.40772e-10, 1.409767e-10, 1.41558e-10, 1.420818e-10, 
    1.426529e-10, 1.427926e-10, 1.4346e-10, 1.429168e-10, 1.438132e-10, 
    1.430511e-10, 1.443703e-10, 1.419999e-10, 1.430287e-10, 1.411649e-10, 
    1.413657e-10, 1.417288e-10, 1.425618e-10, 1.421121e-10, 1.42638e-10, 
    1.414765e-10, 1.408739e-10, 1.40718e-10, 1.404271e-10, 1.407247e-10, 
    1.407005e-10, 1.409852e-10, 1.408937e-10, 1.415773e-10, 1.412101e-10, 
    1.422532e-10, 1.426338e-10, 1.437088e-10, 1.443678e-10, 1.450386e-10, 
    1.453348e-10, 1.454249e-10, 1.454626e-10 ;

 SOIL1N_vr =
  2.497417, 2.49741, 2.497412, 2.497406, 2.497409, 2.497406, 2.497416, 
    2.49741, 2.497414, 2.497416, 2.497396, 2.497406, 2.497385, 2.497391, 
    2.497375, 2.497386, 2.497373, 2.497375, 2.497368, 2.49737, 2.49736, 
    2.497367, 2.497355, 2.497362, 2.497361, 2.497367, 2.497404, 2.497397, 
    2.497404, 2.497403, 2.497404, 2.497409, 2.497412, 2.497418, 2.497416, 
    2.497412, 2.497403, 2.497406, 2.497398, 2.497398, 2.497389, 2.497393, 
    2.497378, 2.497382, 2.49737, 2.497373, 2.49737, 2.497371, 2.49737, 
    2.497375, 2.497373, 2.497377, 2.497392, 2.497388, 2.497402, 2.49741, 
    2.497416, 2.497419, 2.497419, 2.497418, 2.497412, 2.497407, 2.497403, 
    2.497401, 2.497398, 2.497391, 2.497386, 2.497377, 2.497379, 2.497376, 
    2.497373, 2.497369, 2.49737, 2.497368, 2.497376, 2.49737, 2.49738, 
    2.497377, 2.497397, 2.497405, 2.497408, 2.497411, 2.497418, 2.497414, 
    2.497416, 2.497411, 2.497408, 2.49741, 2.497401, 2.497404, 2.497386, 
    2.497394, 2.497374, 2.497379, 2.497373, 2.497375, 2.49737, 2.497375, 
    2.497367, 2.497365, 2.497366, 2.497362, 2.497375, 2.49737, 2.49741, 
    2.497409, 2.497408, 2.497413, 2.497413, 2.497418, 2.497414, 2.497412, 
    2.497408, 2.497405, 2.497403, 2.497398, 2.497392, 2.497384, 2.497378, 
    2.497374, 2.497377, 2.497375, 2.497377, 2.497378, 2.497366, 2.497373, 
    2.497362, 2.497363, 2.497368, 2.497363, 2.497409, 2.497411, 2.497415, 
    2.497411, 2.497418, 2.497414, 2.497412, 2.497404, 2.497402, 2.497401, 
    2.497397, 2.497393, 2.497386, 2.497379, 2.497373, 2.497374, 2.497374, 
    2.497372, 2.497375, 2.497372, 2.497371, 2.497373, 2.497363, 2.497366, 
    2.497363, 2.497365, 2.49741, 2.497408, 2.497409, 2.497407, 2.497408, 
    2.497401, 2.497399, 2.497389, 2.497393, 2.497386, 2.497392, 2.497391, 
    2.497386, 2.497392, 2.49738, 2.497388, 2.497372, 2.497381, 2.497372, 
    2.497373, 2.49737, 2.497368, 2.497365, 2.497359, 2.497361, 2.497356, 
    2.497404, 2.497401, 2.497402, 2.497399, 2.497396, 2.497391, 2.497384, 
    2.497387, 2.497381, 2.49738, 2.497388, 2.497383, 2.4974, 2.497397, 
    2.497398, 2.497404, 2.497386, 2.497395, 2.497378, 2.497383, 2.497368, 
    2.497376, 2.497361, 2.497355, 2.49735, 2.497343, 2.4974, 2.497402, 
    2.497398, 2.497393, 2.497389, 2.497383, 2.497382, 2.497381, 2.497378, 
    2.497376, 2.497381, 2.497375, 2.497396, 2.497385, 2.497403, 2.497397, 
    2.497394, 2.497395, 2.497387, 2.497385, 2.497377, 2.497381, 2.497357, 
    2.497368, 2.497338, 2.497346, 2.497403, 2.4974, 2.497391, 2.497395, 
    2.497382, 2.497379, 2.497377, 2.497374, 2.497373, 2.497371, 2.497375, 
    2.497371, 2.497383, 2.497378, 2.497392, 2.497388, 2.49739, 2.497391, 
    2.497386, 2.497381, 2.49738, 2.497379, 2.497374, 2.497382, 2.497355, 
    2.497372, 2.497397, 2.497392, 2.497391, 2.497393, 2.49738, 2.497385, 
    2.497371, 2.497375, 2.497369, 2.497372, 2.497372, 2.497376, 2.497378, 
    2.497384, 2.497389, 2.497393, 2.497392, 2.497388, 2.49738, 2.497373, 
    2.497375, 2.49737, 2.497383, 2.497378, 2.49738, 2.497374, 2.497387, 
    2.497376, 2.49739, 2.497388, 2.497385, 2.497377, 2.497375, 2.497374, 
    2.497375, 2.49738, 2.497381, 2.497385, 2.497386, 2.497389, 2.497391, 
    2.497389, 2.497386, 2.49738, 2.497374, 2.497368, 2.497366, 2.497359, 
    2.497365, 2.497355, 2.497364, 2.497349, 2.497375, 2.497364, 2.497385, 
    2.497382, 2.497378, 2.497369, 2.497374, 2.497368, 2.497381, 2.497388, 
    2.497389, 2.497393, 2.497389, 2.49739, 2.497386, 2.497387, 2.49738, 
    2.497384, 2.497372, 2.497368, 2.497356, 2.497349, 2.497342, 2.497339, 
    2.497338, 2.497337,
  2.497626, 2.497617, 2.497618, 2.497611, 2.497615, 2.497611, 2.497624, 
    2.497617, 2.497621, 2.497625, 2.497597, 2.497611, 2.497583, 2.497592, 
    2.497571, 2.497585, 2.497567, 2.497571, 2.497561, 2.497564, 2.497551, 
    2.49756, 2.497545, 2.497553, 2.497552, 2.49756, 2.497608, 2.497599, 
    2.497609, 2.497607, 2.497608, 2.497615, 2.497619, 2.497626, 2.497625, 
    2.497619, 2.497607, 2.497611, 2.497601, 2.497601, 2.497589, 2.497594, 
    2.497574, 2.49758, 2.497564, 2.497568, 2.497564, 2.497565, 2.497564, 
    2.49757, 2.497567, 2.497572, 2.497593, 2.497587, 2.497605, 2.497616, 
    2.497623, 2.497629, 2.497628, 2.497627, 2.497619, 2.497613, 2.497608, 
    2.497604, 2.497601, 2.497591, 2.497585, 2.497573, 2.497575, 2.497572, 
    2.497568, 2.497562, 2.497563, 2.497561, 2.497572, 2.497564, 2.497576, 
    2.497573, 2.4976, 2.49761, 2.497614, 2.497618, 2.497627, 2.497621, 
    2.497624, 2.497617, 2.497614, 2.497616, 2.497604, 2.497609, 2.497585, 
    2.497595, 2.497569, 2.497575, 2.497567, 2.497571, 2.497564, 2.49757, 
    2.49756, 2.497557, 2.497559, 2.497553, 2.497571, 2.497564, 2.497616, 
    2.497615, 2.497614, 2.49762, 2.497621, 2.497626, 2.497621, 2.497619, 
    2.497614, 2.49761, 2.497607, 2.4976, 2.497593, 2.497582, 2.497575, 
    2.497569, 2.497572, 2.49757, 2.497573, 2.497574, 2.497558, 2.497567, 
    2.497554, 2.497554, 2.497561, 2.497554, 2.497615, 2.497617, 2.497623, 
    2.497618, 2.497627, 2.497622, 2.497619, 2.497608, 2.497606, 2.497604, 
    2.4976, 2.497594, 2.497584, 2.497576, 2.497568, 2.497569, 2.497568, 
    2.497566, 2.497571, 2.497566, 2.497565, 2.497567, 2.497555, 2.497558, 
    2.497554, 2.497557, 2.497616, 2.497613, 2.497615, 2.497612, 2.497614, 
    2.497605, 2.497602, 2.497589, 2.497594, 2.497586, 2.497593, 2.497592, 
    2.497585, 2.497593, 2.497576, 2.497587, 2.497566, 2.497578, 2.497566, 
    2.497568, 2.497564, 2.497561, 2.497557, 2.49755, 2.497551, 2.497545, 
    2.497609, 2.497605, 2.497606, 2.497602, 2.497598, 2.497592, 2.497582, 
    2.497586, 2.497579, 2.497577, 2.497588, 2.497581, 2.497603, 2.497599, 
    2.497601, 2.497609, 2.497585, 2.497597, 2.497574, 2.497581, 2.497562, 
    2.497571, 2.497552, 2.497544, 2.497537, 2.497528, 2.497603, 2.497606, 
    2.497601, 2.497595, 2.497589, 2.497581, 2.49758, 2.497578, 2.497574, 
    2.497571, 2.497578, 2.49757, 2.497598, 2.497584, 2.497607, 2.4976, 
    2.497595, 2.497597, 2.497586, 2.497583, 2.497573, 2.497578, 2.497546, 
    2.497561, 2.497521, 2.497532, 2.497607, 2.497603, 2.497591, 2.497597, 
    2.49758, 2.497576, 2.497573, 2.497568, 2.497568, 2.497566, 2.49757, 
    2.497566, 2.497581, 2.497574, 2.497592, 2.497588, 2.49759, 2.497592, 
    2.497585, 2.497578, 2.497578, 2.497575, 2.497568, 2.49758, 2.497545, 
    2.497566, 2.497599, 2.497592, 2.497591, 2.497594, 2.497576, 2.497583, 
    2.497566, 2.49757, 2.497562, 2.497566, 2.497567, 2.497572, 2.497575, 
    2.497582, 2.497589, 2.497594, 2.497593, 2.497587, 2.497577, 2.497568, 
    2.49757, 2.497563, 2.497581, 2.497574, 2.497576, 2.497569, 2.497586, 
    2.497571, 2.497589, 2.497588, 2.497583, 2.497573, 2.497571, 2.497569, 
    2.49757, 2.497577, 2.497578, 2.497583, 2.497584, 2.497588, 2.497591, 
    2.497588, 2.497586, 2.497577, 2.497569, 2.497561, 2.497559, 2.497549, 
    2.497557, 2.497544, 2.497555, 2.497536, 2.497571, 2.497556, 2.497583, 
    2.49758, 2.497575, 2.497562, 2.497569, 2.497561, 2.497578, 2.497587, 
    2.497589, 2.497593, 2.497589, 2.49759, 2.497585, 2.497587, 2.497577, 
    2.497582, 2.497567, 2.497561, 2.497546, 2.497536, 2.497527, 2.497522, 
    2.497521, 2.49752,
  2.497841, 2.497832, 2.497833, 2.497826, 2.49783, 2.497825, 2.497839, 
    2.497831, 2.497836, 2.49784, 2.497811, 2.497825, 2.497796, 2.497805, 
    2.497782, 2.497797, 2.497779, 2.497782, 2.497772, 2.497775, 2.497761, 
    2.49777, 2.497754, 2.497763, 2.497762, 2.497771, 2.497823, 2.497813, 
    2.497823, 2.497822, 2.497822, 2.49783, 2.497834, 2.497842, 2.49784, 
    2.497834, 2.497821, 2.497826, 2.497814, 2.497814, 2.497802, 2.497808, 
    2.497786, 2.497792, 2.497775, 2.497779, 2.497775, 2.497776, 2.497775, 
    2.497781, 2.497779, 2.497784, 2.497806, 2.4978, 2.497819, 2.497831, 
    2.497839, 2.497844, 2.497844, 2.497842, 2.497834, 2.497827, 2.497822, 
    2.497818, 2.497814, 2.497803, 2.497798, 2.497785, 2.497787, 2.497783, 
    2.49778, 2.497773, 2.497774, 2.497772, 2.497783, 2.497776, 2.497789, 
    2.497785, 2.497813, 2.497824, 2.497829, 2.497833, 2.497843, 2.497836, 
    2.497839, 2.497832, 2.497828, 2.49783, 2.497818, 2.497823, 2.497797, 
    2.497808, 2.49778, 2.497787, 2.497778, 2.497783, 2.497775, 2.497782, 
    2.497771, 2.497768, 2.49777, 2.497763, 2.497782, 2.497775, 2.49783, 
    2.49783, 2.497828, 2.497835, 2.497836, 2.497842, 2.497836, 2.497834, 
    2.497828, 2.497825, 2.497821, 2.497814, 2.497806, 2.497794, 2.497786, 
    2.497781, 2.497784, 2.497781, 2.497785, 2.497786, 2.497769, 2.497779, 
    2.497764, 2.497765, 2.497772, 2.497765, 2.49783, 2.497832, 2.497838, 
    2.497833, 2.497843, 2.497837, 2.497834, 2.497823, 2.49782, 2.497818, 
    2.497813, 2.497807, 2.497797, 2.497788, 2.497779, 2.49778, 2.49778, 
    2.497778, 2.497782, 2.497777, 2.497776, 2.497779, 2.497765, 2.497769, 
    2.497765, 2.497767, 2.497831, 2.497828, 2.49783, 2.497826, 2.497829, 
    2.497819, 2.497816, 2.497802, 2.497807, 2.497798, 2.497806, 2.497805, 
    2.497798, 2.497806, 2.497788, 2.4978, 2.497778, 2.49779, 2.497777, 
    2.497779, 2.497776, 2.497772, 2.497768, 2.49776, 2.497762, 2.497755, 
    2.497823, 2.497819, 2.497819, 2.497815, 2.497812, 2.497805, 2.497794, 
    2.497798, 2.497791, 2.497789, 2.497801, 2.497794, 2.497816, 2.497813, 
    2.497815, 2.497823, 2.497797, 2.49781, 2.497786, 2.497793, 2.497773, 
    2.497783, 2.497763, 2.497754, 2.497746, 2.497736, 2.497817, 2.49782, 
    2.497815, 2.497808, 2.497801, 2.497793, 2.497792, 2.49779, 2.497786, 
    2.497783, 2.49779, 2.497782, 2.497812, 2.497796, 2.497821, 2.497813, 
    2.497808, 2.49781, 2.497799, 2.497796, 2.497785, 2.497791, 2.497756, 
    2.497771, 2.497729, 2.497741, 2.497821, 2.497817, 2.497804, 2.49781, 
    2.497792, 2.497788, 2.497784, 2.49778, 2.497779, 2.497777, 2.497781, 
    2.497777, 2.497793, 2.497786, 2.497805, 2.497801, 2.497803, 2.497805, 
    2.497798, 2.49779, 2.49779, 2.497787, 2.49778, 2.497792, 2.497754, 
    2.497778, 2.497813, 2.497806, 2.497805, 2.497807, 2.497788, 2.497795, 
    2.497777, 2.497782, 2.497774, 2.497778, 2.497778, 2.497783, 2.497787, 
    2.497795, 2.497802, 2.497807, 2.497806, 2.4978, 2.497789, 2.497779, 
    2.497782, 2.497774, 2.497794, 2.497785, 2.497789, 2.49778, 2.497798, 
    2.497783, 2.497802, 2.497801, 2.497795, 2.497785, 2.497782, 2.49778, 
    2.497782, 2.497789, 2.49779, 2.497796, 2.497797, 2.497801, 2.497804, 
    2.497801, 2.497798, 2.497789, 2.497781, 2.497772, 2.49777, 2.49776, 
    2.497768, 2.497754, 2.497766, 2.497746, 2.497782, 2.497766, 2.497795, 
    2.497792, 2.497786, 2.497773, 2.49778, 2.497772, 2.49779, 2.4978, 
    2.497802, 2.497807, 2.497802, 2.497802, 2.497798, 2.497799, 2.497789, 
    2.497794, 2.497778, 2.497772, 2.497756, 2.497746, 2.497735, 2.49773, 
    2.497729, 2.497729,
  2.498013, 2.498003, 2.498005, 2.497998, 2.498002, 2.497997, 2.498011, 
    2.498003, 2.498008, 2.498012, 2.497983, 2.497997, 2.497968, 2.497977, 
    2.497954, 2.49797, 2.497951, 2.497955, 2.497944, 2.497947, 2.497934, 
    2.497943, 2.497927, 2.497936, 2.497934, 2.497943, 2.497994, 2.497985, 
    2.497995, 2.497994, 2.497994, 2.498002, 2.498006, 2.498013, 2.498012, 
    2.498006, 2.497993, 2.497998, 2.497986, 2.497987, 2.497974, 2.49798, 
    2.497958, 2.497964, 2.497947, 2.497952, 2.497947, 2.497948, 2.497947, 
    2.497954, 2.497951, 2.497957, 2.497978, 2.497972, 2.497991, 2.498003, 
    2.498011, 2.498016, 2.498015, 2.498014, 2.498006, 2.497999, 2.497994, 
    2.49799, 2.497987, 2.497976, 2.49797, 2.497957, 2.49796, 2.497956, 
    2.497952, 2.497946, 2.497947, 2.497944, 2.497956, 2.497948, 2.497961, 
    2.497957, 2.497986, 2.497996, 2.498001, 2.498005, 2.498015, 2.498008, 
    2.498011, 2.498004, 2.498, 2.498002, 2.49799, 2.497995, 2.49797, 2.49798, 
    2.497952, 2.497959, 2.497951, 2.497955, 2.497948, 2.497954, 2.497943, 
    2.49794, 2.497942, 2.497936, 2.497955, 2.497947, 2.498002, 2.498002, 
    2.498, 2.498007, 2.498008, 2.498013, 2.498008, 2.498006, 2.498, 2.497997, 
    2.497993, 2.497986, 2.497978, 2.497967, 2.497959, 2.497953, 2.497957, 
    2.497954, 2.497957, 2.497958, 2.497941, 2.497951, 2.497936, 2.497937, 
    2.497944, 2.497937, 2.498002, 2.498003, 2.49801, 2.498005, 2.498014, 
    2.498009, 2.498006, 2.497995, 2.497992, 2.49799, 2.497985, 2.497979, 
    2.497969, 2.49796, 2.497952, 2.497952, 2.497952, 2.49795, 2.497955, 
    2.497949, 2.497949, 2.497951, 2.497937, 2.497941, 2.497937, 2.49794, 
    2.498003, 2.498, 2.498002, 2.497998, 2.498001, 2.497991, 2.497988, 
    2.497974, 2.497979, 2.49797, 2.497978, 2.497977, 2.49797, 2.497978, 
    2.49796, 2.497972, 2.49795, 2.497962, 2.497949, 2.497952, 2.497948, 
    2.497944, 2.49794, 2.497932, 2.497934, 2.497927, 2.497995, 2.497991, 
    2.497992, 2.497987, 2.497984, 2.497977, 2.497966, 2.49797, 2.497963, 
    2.497961, 2.497973, 2.497966, 2.497988, 2.497985, 2.497987, 2.497995, 
    2.497969, 2.497983, 2.497958, 2.497966, 2.497945, 2.497955, 2.497935, 
    2.497926, 2.497918, 2.497909, 2.497989, 2.497992, 2.497987, 2.49798, 
    2.497973, 2.497965, 2.497964, 2.497963, 2.497959, 2.497955, 2.497962, 
    2.497954, 2.497984, 2.497968, 2.497993, 2.497985, 2.49798, 2.497983, 
    2.497971, 2.497968, 2.497957, 2.497963, 2.497929, 2.497944, 2.497902, 
    2.497914, 2.497993, 2.497989, 2.497976, 2.497982, 2.497965, 2.49796, 
    2.497957, 2.497952, 2.497952, 2.497949, 2.497953, 2.497949, 2.497965, 
    2.497958, 2.497977, 2.497973, 2.497975, 2.497977, 2.49797, 2.497962, 
    2.497962, 2.497959, 2.497952, 2.497964, 2.497927, 2.49795, 2.497985, 
    2.497978, 2.497977, 2.497979, 2.497961, 2.497967, 2.497949, 2.497954, 
    2.497946, 2.49795, 2.497951, 2.497956, 2.497959, 2.497967, 2.497974, 
    2.497979, 2.497978, 2.497972, 2.497962, 2.497952, 2.497954, 2.497947, 
    2.497966, 2.497958, 2.497961, 2.497953, 2.497971, 2.497955, 2.497974, 
    2.497973, 2.497967, 2.497957, 2.497955, 2.497952, 2.497954, 2.497961, 
    2.497962, 2.497968, 2.497969, 2.497973, 2.497976, 2.497973, 2.49797, 
    2.497961, 2.497953, 2.497944, 2.497942, 2.497932, 2.49794, 2.497926, 
    2.497938, 2.497918, 2.497954, 2.497939, 2.497967, 2.497964, 2.497959, 
    2.497946, 2.497953, 2.497945, 2.497962, 2.497972, 2.497974, 2.497979, 
    2.497974, 2.497974, 2.49797, 2.497972, 2.497961, 2.497967, 2.497951, 
    2.497945, 2.497928, 2.497918, 2.497908, 2.497903, 2.497902, 2.497901,
  2.498213, 2.498205, 2.498207, 2.4982, 2.498204, 2.498199, 2.498212, 
    2.498205, 2.498209, 2.498213, 2.498187, 2.498199, 2.498174, 2.498182, 
    2.498161, 2.498175, 2.498159, 2.498162, 2.498152, 2.498155, 2.498143, 
    2.498151, 2.498137, 2.498145, 2.498144, 2.498151, 2.498197, 2.498188, 
    2.498198, 2.498196, 2.498197, 2.498204, 2.498207, 2.498214, 2.498213, 
    2.498207, 2.498196, 2.4982, 2.49819, 2.49819, 2.498179, 2.498184, 
    2.498165, 2.49817, 2.498155, 2.498159, 2.498155, 2.498156, 2.498155, 
    2.498161, 2.498158, 2.498163, 2.498183, 2.498177, 2.498194, 2.498204, 
    2.498211, 2.498216, 2.498215, 2.498214, 2.498207, 2.498201, 2.498196, 
    2.498193, 2.49819, 2.49818, 2.498175, 2.498164, 2.498166, 2.498163, 
    2.498159, 2.498154, 2.498154, 2.498152, 2.498163, 2.498156, 2.498167, 
    2.498164, 2.498189, 2.498199, 2.498203, 2.498206, 2.498215, 2.498209, 
    2.498211, 2.498206, 2.498202, 2.498204, 2.498193, 2.498197, 2.498175, 
    2.498185, 2.49816, 2.498166, 2.498158, 2.498162, 2.498155, 2.498161, 
    2.498151, 2.498149, 2.49815, 2.498145, 2.498162, 2.498155, 2.498204, 
    2.498204, 2.498202, 2.498208, 2.498209, 2.498214, 2.498209, 2.498207, 
    2.498202, 2.498199, 2.498196, 2.498189, 2.498182, 2.498172, 2.498165, 
    2.49816, 2.498163, 2.498161, 2.498164, 2.498165, 2.49815, 2.498158, 
    2.498145, 2.498146, 2.498152, 2.498146, 2.498204, 2.498205, 2.498211, 
    2.498206, 2.498214, 2.49821, 2.498207, 2.498197, 2.498195, 2.498193, 
    2.498189, 2.498183, 2.498174, 2.498166, 2.498159, 2.498159, 2.498159, 
    2.498158, 2.498162, 2.498157, 2.498156, 2.498158, 2.498146, 2.49815, 
    2.498146, 2.498148, 2.498204, 2.498202, 2.498203, 2.4982, 2.498202, 
    2.498194, 2.498191, 2.498178, 2.498184, 2.498175, 2.498183, 2.498182, 
    2.498175, 2.498182, 2.498167, 2.498177, 2.498158, 2.498168, 2.498157, 
    2.498159, 2.498156, 2.498152, 2.498149, 2.498142, 2.498143, 2.498137, 
    2.498198, 2.498194, 2.498194, 2.498191, 2.498188, 2.498182, 2.498172, 
    2.498176, 2.498169, 2.498168, 2.498178, 2.498172, 2.498192, 2.498188, 
    2.49819, 2.498197, 2.498175, 2.498186, 2.498165, 2.498171, 2.498153, 
    2.498162, 2.498144, 2.498137, 2.498129, 2.498121, 2.498192, 2.498194, 
    2.49819, 2.498184, 2.498178, 2.498171, 2.49817, 2.498169, 2.498165, 
    2.498162, 2.498168, 2.498161, 2.498188, 2.498174, 2.498195, 2.498189, 
    2.498184, 2.498186, 2.498176, 2.498174, 2.498164, 2.498169, 2.498138, 
    2.498152, 2.498115, 2.498125, 2.498195, 2.498192, 2.498181, 2.498186, 
    2.49817, 2.498167, 2.498163, 2.498159, 2.498159, 2.498157, 2.498161, 
    2.498157, 2.498171, 2.498165, 2.498182, 2.498178, 2.49818, 2.498182, 
    2.498175, 2.498168, 2.498168, 2.498166, 2.498159, 2.49817, 2.498137, 
    2.498158, 2.498188, 2.498182, 2.498181, 2.498184, 2.498167, 2.498173, 
    2.498157, 2.498161, 2.498154, 2.498158, 2.498158, 2.498163, 2.498165, 
    2.498173, 2.498179, 2.498183, 2.498182, 2.498177, 2.498168, 2.498159, 
    2.498161, 2.498154, 2.498172, 2.498164, 2.498167, 2.49816, 2.498176, 
    2.498162, 2.498179, 2.498178, 2.498173, 2.498164, 2.498162, 2.49816, 
    2.498161, 2.498168, 2.498169, 2.498173, 2.498174, 2.498178, 2.498181, 
    2.498178, 2.498175, 2.498168, 2.49816, 2.498152, 2.498151, 2.498142, 
    2.498149, 2.498137, 2.498147, 2.498129, 2.498162, 2.498147, 2.498173, 
    2.49817, 2.498165, 2.498154, 2.49816, 2.498153, 2.498169, 2.498177, 
    2.498179, 2.498183, 2.498179, 2.498179, 2.498175, 2.498177, 2.498167, 
    2.498172, 2.498158, 2.498153, 2.498138, 2.498129, 2.49812, 2.498116, 
    2.498114, 2.498114,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1_HR_S2 =
  6.139198e-08, 6.166193e-08, 6.160945e-08, 6.182718e-08, 6.170639e-08, 
    6.184897e-08, 6.144671e-08, 6.167265e-08, 6.152841e-08, 6.141628e-08, 
    6.224973e-08, 6.183689e-08, 6.267852e-08, 6.241524e-08, 6.307661e-08, 
    6.263755e-08, 6.316512e-08, 6.306393e-08, 6.33685e-08, 6.328124e-08, 
    6.367082e-08, 6.340877e-08, 6.387275e-08, 6.360823e-08, 6.364962e-08, 
    6.340012e-08, 6.191997e-08, 6.219834e-08, 6.190348e-08, 6.194317e-08, 
    6.192536e-08, 6.17089e-08, 6.159981e-08, 6.137134e-08, 6.141282e-08, 
    6.158062e-08, 6.196102e-08, 6.183189e-08, 6.215732e-08, 6.214997e-08, 
    6.251226e-08, 6.234892e-08, 6.295784e-08, 6.278477e-08, 6.328489e-08, 
    6.315911e-08, 6.327897e-08, 6.324263e-08, 6.327945e-08, 6.309499e-08, 
    6.317403e-08, 6.301171e-08, 6.237951e-08, 6.256531e-08, 6.201116e-08, 
    6.167795e-08, 6.145662e-08, 6.129956e-08, 6.132176e-08, 6.136409e-08, 
    6.15816e-08, 6.17861e-08, 6.194195e-08, 6.20462e-08, 6.214891e-08, 
    6.245984e-08, 6.262439e-08, 6.299284e-08, 6.292634e-08, 6.303899e-08, 
    6.31466e-08, 6.332728e-08, 6.329753e-08, 6.337714e-08, 6.303601e-08, 
    6.326273e-08, 6.288847e-08, 6.299083e-08, 6.217687e-08, 6.186672e-08, 
    6.173492e-08, 6.161954e-08, 6.133883e-08, 6.153268e-08, 6.145627e-08, 
    6.163806e-08, 6.175357e-08, 6.169644e-08, 6.204905e-08, 6.191197e-08, 
    6.263414e-08, 6.232308e-08, 6.313405e-08, 6.293999e-08, 6.318056e-08, 
    6.30578e-08, 6.326815e-08, 6.307884e-08, 6.340677e-08, 6.347817e-08, 
    6.342938e-08, 6.361681e-08, 6.306834e-08, 6.327898e-08, 6.169484e-08, 
    6.170416e-08, 6.174757e-08, 6.155675e-08, 6.154508e-08, 6.137021e-08, 
    6.152581e-08, 6.159207e-08, 6.176027e-08, 6.185977e-08, 6.195435e-08, 
    6.216229e-08, 6.239453e-08, 6.271927e-08, 6.295257e-08, 6.310896e-08, 
    6.301306e-08, 6.309772e-08, 6.300308e-08, 6.295872e-08, 6.345142e-08, 
    6.317477e-08, 6.358985e-08, 6.356689e-08, 6.337903e-08, 6.356947e-08, 
    6.171071e-08, 6.165708e-08, 6.147091e-08, 6.161661e-08, 6.135116e-08, 
    6.149975e-08, 6.158519e-08, 6.191484e-08, 6.198726e-08, 6.205442e-08, 
    6.218706e-08, 6.235727e-08, 6.265589e-08, 6.291569e-08, 6.315286e-08, 
    6.313548e-08, 6.31416e-08, 6.319458e-08, 6.306335e-08, 6.321613e-08, 
    6.324178e-08, 6.317473e-08, 6.356381e-08, 6.345265e-08, 6.35664e-08, 
    6.349402e-08, 6.167451e-08, 6.176474e-08, 6.171599e-08, 6.180766e-08, 
    6.174308e-08, 6.203027e-08, 6.211638e-08, 6.251928e-08, 6.235393e-08, 
    6.261709e-08, 6.238066e-08, 6.242255e-08, 6.262568e-08, 6.239343e-08, 
    6.290137e-08, 6.255701e-08, 6.319664e-08, 6.285278e-08, 6.32182e-08, 
    6.315184e-08, 6.32617e-08, 6.33601e-08, 6.348389e-08, 6.371231e-08, 
    6.365941e-08, 6.385043e-08, 6.189924e-08, 6.201627e-08, 6.200596e-08, 
    6.212843e-08, 6.2219e-08, 6.24153e-08, 6.273014e-08, 6.261175e-08, 
    6.28291e-08, 6.287274e-08, 6.254253e-08, 6.274527e-08, 6.209459e-08, 
    6.219972e-08, 6.213713e-08, 6.190847e-08, 6.263904e-08, 6.226412e-08, 
    6.295642e-08, 6.275332e-08, 6.334607e-08, 6.30513e-08, 6.36303e-08, 
    6.387783e-08, 6.411076e-08, 6.438301e-08, 6.208013e-08, 6.200062e-08, 
    6.214299e-08, 6.233998e-08, 6.252274e-08, 6.276571e-08, 6.279057e-08, 
    6.283609e-08, 6.295399e-08, 6.305312e-08, 6.285049e-08, 6.307798e-08, 
    6.222412e-08, 6.267158e-08, 6.197056e-08, 6.218166e-08, 6.232837e-08, 
    6.226401e-08, 6.259822e-08, 6.267699e-08, 6.299708e-08, 6.283161e-08, 
    6.381674e-08, 6.33809e-08, 6.459028e-08, 6.425232e-08, 6.197283e-08, 
    6.207986e-08, 6.245234e-08, 6.227511e-08, 6.278193e-08, 6.290668e-08, 
    6.300809e-08, 6.313773e-08, 6.315172e-08, 6.322854e-08, 6.310267e-08, 
    6.322357e-08, 6.276623e-08, 6.29706e-08, 6.240975e-08, 6.254626e-08, 
    6.248347e-08, 6.241458e-08, 6.262718e-08, 6.285368e-08, 6.285851e-08, 
    6.293114e-08, 6.313581e-08, 6.278398e-08, 6.387301e-08, 6.320047e-08, 
    6.219656e-08, 6.240271e-08, 6.243215e-08, 6.235229e-08, 6.289418e-08, 
    6.269784e-08, 6.322666e-08, 6.308374e-08, 6.331792e-08, 6.320155e-08, 
    6.318443e-08, 6.303497e-08, 6.294192e-08, 6.270684e-08, 6.251556e-08, 
    6.236387e-08, 6.239915e-08, 6.256577e-08, 6.286754e-08, 6.3153e-08, 
    6.309047e-08, 6.330012e-08, 6.274518e-08, 6.297788e-08, 6.288795e-08, 
    6.312245e-08, 6.260861e-08, 6.30462e-08, 6.249675e-08, 6.254493e-08, 
    6.269394e-08, 6.299367e-08, 6.305997e-08, 6.313078e-08, 6.308709e-08, 
    6.287519e-08, 6.284047e-08, 6.269031e-08, 6.264886e-08, 6.253444e-08, 
    6.243971e-08, 6.252626e-08, 6.261715e-08, 6.287528e-08, 6.310789e-08, 
    6.33615e-08, 6.342356e-08, 6.37199e-08, 6.347868e-08, 6.387675e-08, 
    6.353834e-08, 6.412414e-08, 6.307155e-08, 6.352837e-08, 6.270071e-08, 
    6.278988e-08, 6.295116e-08, 6.332105e-08, 6.312135e-08, 6.335489e-08, 
    6.283911e-08, 6.257152e-08, 6.250227e-08, 6.23731e-08, 6.250523e-08, 
    6.249448e-08, 6.262091e-08, 6.258028e-08, 6.288385e-08, 6.272079e-08, 
    6.3184e-08, 6.335304e-08, 6.383041e-08, 6.412306e-08, 6.442093e-08, 
    6.455244e-08, 6.459247e-08, 6.46092e-08 ;

 SOIL1_HR_S3 =
  7.285347e-10, 7.317394e-10, 7.311164e-10, 7.337012e-10, 7.322674e-10, 
    7.339599e-10, 7.291844e-10, 7.318667e-10, 7.301544e-10, 7.288232e-10, 
    7.387176e-10, 7.338165e-10, 7.438081e-10, 7.406825e-10, 7.485342e-10, 
    7.433218e-10, 7.495852e-10, 7.483837e-10, 7.519997e-10, 7.509637e-10, 
    7.55589e-10, 7.524777e-10, 7.579865e-10, 7.548459e-10, 7.553372e-10, 
    7.523752e-10, 7.348028e-10, 7.381075e-10, 7.34607e-10, 7.350782e-10, 
    7.348668e-10, 7.32297e-10, 7.31002e-10, 7.282898e-10, 7.287821e-10, 
    7.307742e-10, 7.352901e-10, 7.337571e-10, 7.376205e-10, 7.375333e-10, 
    7.418344e-10, 7.398951e-10, 7.471243e-10, 7.450696e-10, 7.51007e-10, 
    7.495138e-10, 7.509369e-10, 7.505053e-10, 7.509425e-10, 7.487526e-10, 
    7.496908e-10, 7.477638e-10, 7.402583e-10, 7.424641e-10, 7.358853e-10, 
    7.319297e-10, 7.293021e-10, 7.274376e-10, 7.277012e-10, 7.282037e-10, 
    7.307859e-10, 7.332136e-10, 7.350637e-10, 7.363013e-10, 7.375207e-10, 
    7.41212e-10, 7.431655e-10, 7.475398e-10, 7.467503e-10, 7.480877e-10, 
    7.493652e-10, 7.515103e-10, 7.511572e-10, 7.521023e-10, 7.480523e-10, 
    7.50744e-10, 7.463006e-10, 7.475159e-10, 7.378526e-10, 7.341707e-10, 
    7.32606e-10, 7.312362e-10, 7.279038e-10, 7.302051e-10, 7.292979e-10, 
    7.314561e-10, 7.328274e-10, 7.321492e-10, 7.363352e-10, 7.347077e-10, 
    7.432813e-10, 7.395884e-10, 7.492162e-10, 7.469123e-10, 7.497685e-10, 
    7.48311e-10, 7.508082e-10, 7.485608e-10, 7.52454e-10, 7.533018e-10, 
    7.527224e-10, 7.549478e-10, 7.484362e-10, 7.509369e-10, 7.321302e-10, 
    7.322408e-10, 7.327561e-10, 7.304908e-10, 7.303523e-10, 7.282763e-10, 
    7.301235e-10, 7.309101e-10, 7.329069e-10, 7.340881e-10, 7.352108e-10, 
    7.376796e-10, 7.404367e-10, 7.44292e-10, 7.470617e-10, 7.489183e-10, 
    7.477798e-10, 7.487849e-10, 7.476613e-10, 7.471347e-10, 7.529841e-10, 
    7.496996e-10, 7.546277e-10, 7.54355e-10, 7.521248e-10, 7.543857e-10, 
    7.323185e-10, 7.316819e-10, 7.294718e-10, 7.312014e-10, 7.280502e-10, 
    7.298141e-10, 7.308284e-10, 7.347418e-10, 7.356016e-10, 7.363989e-10, 
    7.379735e-10, 7.399943e-10, 7.435394e-10, 7.466239e-10, 7.494396e-10, 
    7.492332e-10, 7.493059e-10, 7.499349e-10, 7.483768e-10, 7.501907e-10, 
    7.504952e-10, 7.496992e-10, 7.543184e-10, 7.529988e-10, 7.543492e-10, 
    7.534899e-10, 7.318888e-10, 7.329599e-10, 7.323812e-10, 7.334695e-10, 
    7.327028e-10, 7.361123e-10, 7.371345e-10, 7.419177e-10, 7.399546e-10, 
    7.430788e-10, 7.402719e-10, 7.407693e-10, 7.431809e-10, 7.404236e-10, 
    7.464538e-10, 7.423657e-10, 7.499594e-10, 7.45877e-10, 7.502152e-10, 
    7.494274e-10, 7.507318e-10, 7.519e-10, 7.533696e-10, 7.560815e-10, 
    7.554535e-10, 7.577213e-10, 7.345567e-10, 7.35946e-10, 7.358236e-10, 
    7.372775e-10, 7.383528e-10, 7.406832e-10, 7.44421e-10, 7.430154e-10, 
    7.455959e-10, 7.461139e-10, 7.421936e-10, 7.446007e-10, 7.368758e-10, 
    7.381239e-10, 7.373808e-10, 7.346663e-10, 7.433394e-10, 7.388884e-10, 
    7.471074e-10, 7.446962e-10, 7.517335e-10, 7.482338e-10, 7.551078e-10, 
    7.580467e-10, 7.608122e-10, 7.640446e-10, 7.367042e-10, 7.357602e-10, 
    7.374504e-10, 7.39789e-10, 7.419587e-10, 7.448433e-10, 7.451384e-10, 
    7.456788e-10, 7.470786e-10, 7.482555e-10, 7.458498e-10, 7.485505e-10, 
    7.384135e-10, 7.437257e-10, 7.354033e-10, 7.379095e-10, 7.396511e-10, 
    7.388871e-10, 7.428548e-10, 7.4379e-10, 7.475902e-10, 7.456256e-10, 
    7.573214e-10, 7.521468e-10, 7.665055e-10, 7.624929e-10, 7.354304e-10, 
    7.367009e-10, 7.411229e-10, 7.390189e-10, 7.450358e-10, 7.465169e-10, 
    7.477208e-10, 7.4926e-10, 7.494261e-10, 7.50338e-10, 7.488437e-10, 
    7.50279e-10, 7.448495e-10, 7.472757e-10, 7.406174e-10, 7.42238e-10, 
    7.414924e-10, 7.406747e-10, 7.431986e-10, 7.458876e-10, 7.45945e-10, 
    7.468072e-10, 7.492372e-10, 7.450602e-10, 7.579894e-10, 7.500048e-10, 
    7.380864e-10, 7.405337e-10, 7.408832e-10, 7.399352e-10, 7.463684e-10, 
    7.440374e-10, 7.503158e-10, 7.486189e-10, 7.513992e-10, 7.500177e-10, 
    7.498144e-10, 7.4804e-10, 7.469353e-10, 7.441444e-10, 7.418735e-10, 
    7.400727e-10, 7.404914e-10, 7.424695e-10, 7.460521e-10, 7.494412e-10, 
    7.486988e-10, 7.511879e-10, 7.445995e-10, 7.473622e-10, 7.462945e-10, 
    7.490785e-10, 7.429781e-10, 7.481733e-10, 7.416502e-10, 7.422221e-10, 
    7.439911e-10, 7.475496e-10, 7.483368e-10, 7.491774e-10, 7.486587e-10, 
    7.46143e-10, 7.457309e-10, 7.439481e-10, 7.43456e-10, 7.420976e-10, 
    7.409731e-10, 7.420005e-10, 7.430796e-10, 7.46144e-10, 7.489057e-10, 
    7.519166e-10, 7.526534e-10, 7.561717e-10, 7.533078e-10, 7.58034e-10, 
    7.540161e-10, 7.609711e-10, 7.484742e-10, 7.538977e-10, 7.440716e-10, 
    7.451302e-10, 7.470449e-10, 7.514363e-10, 7.490654e-10, 7.518381e-10, 
    7.457147e-10, 7.425378e-10, 7.417157e-10, 7.401821e-10, 7.417508e-10, 
    7.416232e-10, 7.431242e-10, 7.426419e-10, 7.462458e-10, 7.443099e-10, 
    7.498093e-10, 7.518162e-10, 7.574837e-10, 7.609582e-10, 7.644948e-10, 
    7.660562e-10, 7.665314e-10, 7.667301e-10 ;

 SOIL2C =
  5.784045, 5.784051, 5.78405, 5.784055, 5.784052, 5.784055, 5.784046, 
    5.784051, 5.784048, 5.784045, 5.784065, 5.784055, 5.784075, 5.784069, 
    5.784084, 5.784074, 5.784086, 5.784084, 5.784091, 5.784089, 5.784098, 
    5.784092, 5.784103, 5.784097, 5.784098, 5.784091, 5.784057, 5.784063, 
    5.784057, 5.784058, 5.784057, 5.784052, 5.78405, 5.784044, 5.784045, 
    5.784049, 5.784058, 5.784055, 5.784062, 5.784062, 5.784071, 5.784067, 
    5.784081, 5.784077, 5.784089, 5.784086, 5.784089, 5.784088, 5.784089, 
    5.784084, 5.784086, 5.784082, 5.784068, 5.784072, 5.784059, 5.784051, 
    5.784046, 5.784042, 5.784043, 5.784044, 5.784049, 5.784054, 5.784058, 
    5.78406, 5.784062, 5.78407, 5.784073, 5.784082, 5.784081, 5.784083, 
    5.784086, 5.78409, 5.784089, 5.784091, 5.784083, 5.784089, 5.78408, 
    5.784082, 5.784063, 5.784056, 5.784052, 5.78405, 5.784043, 5.784048, 
    5.784046, 5.78405, 5.784053, 5.784052, 5.78406, 5.784057, 5.784074, 
    5.784066, 5.784085, 5.784081, 5.784087, 5.784084, 5.784089, 5.784084, 
    5.784092, 5.784093, 5.784092, 5.784097, 5.784084, 5.784089, 5.784051, 
    5.784052, 5.784053, 5.784049, 5.784048, 5.784044, 5.784048, 5.784049, 
    5.784053, 5.784056, 5.784058, 5.784062, 5.784068, 5.784076, 5.784081, 
    5.784085, 5.784082, 5.784084, 5.784082, 5.784081, 5.784093, 5.784086, 
    5.784096, 5.784096, 5.784091, 5.784096, 5.784052, 5.784051, 5.784046, 
    5.78405, 5.784044, 5.784047, 5.784049, 5.784057, 5.784059, 5.78406, 
    5.784063, 5.784067, 5.784074, 5.784081, 5.784086, 5.784085, 5.784086, 
    5.784087, 5.784084, 5.784087, 5.784088, 5.784086, 5.784095, 5.784093, 
    5.784096, 5.784094, 5.784051, 5.784053, 5.784052, 5.784054, 5.784053, 
    5.78406, 5.784061, 5.784071, 5.784067, 5.784073, 5.784068, 5.784069, 
    5.784073, 5.784068, 5.78408, 5.784072, 5.784087, 5.784079, 5.784087, 
    5.784086, 5.784089, 5.784091, 5.784093, 5.784099, 5.784098, 5.784102, 
    5.784057, 5.784059, 5.784059, 5.784062, 5.784064, 5.784069, 5.784076, 
    5.784073, 5.784078, 5.784079, 5.784071, 5.784076, 5.784061, 5.784063, 
    5.784062, 5.784057, 5.784074, 5.784065, 5.784081, 5.784077, 5.784091, 
    5.784083, 5.784097, 5.784103, 5.784108, 5.784115, 5.78406, 5.784059, 
    5.784062, 5.784067, 5.784071, 5.784077, 5.784077, 5.784079, 5.784081, 
    5.784083, 5.784079, 5.784084, 5.784064, 5.784075, 5.784058, 5.784063, 
    5.784067, 5.784065, 5.784073, 5.784075, 5.784082, 5.784078, 5.784101, 
    5.784091, 5.78412, 5.784111, 5.784058, 5.78406, 5.78407, 5.784065, 
    5.784077, 5.78408, 5.784082, 5.784085, 5.784086, 5.784088, 5.784085, 
    5.784088, 5.784077, 5.784081, 5.784069, 5.784071, 5.78407, 5.784069, 
    5.784073, 5.784079, 5.784079, 5.784081, 5.784085, 5.784077, 5.784103, 
    5.784087, 5.784063, 5.784068, 5.784069, 5.784067, 5.78408, 5.784075, 
    5.784088, 5.784084, 5.78409, 5.784087, 5.784087, 5.784083, 5.784081, 
    5.784075, 5.784071, 5.784067, 5.784068, 5.784072, 5.784079, 5.784086, 
    5.784084, 5.784089, 5.784076, 5.784082, 5.78408, 5.784085, 5.784073, 
    5.784083, 5.78407, 5.784071, 5.784075, 5.784082, 5.784084, 5.784085, 
    5.784084, 5.78408, 5.784079, 5.784075, 5.784074, 5.784071, 5.784069, 
    5.784071, 5.784073, 5.78408, 5.784085, 5.784091, 5.784092, 5.784099, 
    5.784093, 5.784103, 5.784095, 5.784109, 5.784084, 5.784095, 5.784075, 
    5.784077, 5.784081, 5.78409, 5.784085, 5.784091, 5.784079, 5.784072, 
    5.78407, 5.784068, 5.78407, 5.78407, 5.784073, 5.784072, 5.78408, 
    5.784076, 5.784087, 5.784091, 5.784101, 5.784109, 5.784116, 5.784119, 
    5.78412, 5.78412 ;

 SOIL2C_TO_SOIL1C =
  1.086144e-09, 1.090923e-09, 1.089994e-09, 1.093849e-09, 1.091711e-09, 
    1.094235e-09, 1.087113e-09, 1.091113e-09, 1.088559e-09, 1.086574e-09, 
    1.101331e-09, 1.094021e-09, 1.108923e-09, 1.104261e-09, 1.115971e-09, 
    1.108197e-09, 1.117538e-09, 1.115746e-09, 1.121139e-09, 1.119594e-09, 
    1.126492e-09, 1.121852e-09, 1.130067e-09, 1.125384e-09, 1.126116e-09, 
    1.121699e-09, 1.095492e-09, 1.100421e-09, 1.0952e-09, 1.095903e-09, 
    1.095588e-09, 1.091755e-09, 1.089824e-09, 1.085778e-09, 1.086513e-09, 
    1.089484e-09, 1.096219e-09, 1.093933e-09, 1.099694e-09, 1.099564e-09, 
    1.105979e-09, 1.103087e-09, 1.113868e-09, 1.110804e-09, 1.119659e-09, 
    1.117432e-09, 1.119554e-09, 1.11891e-09, 1.119562e-09, 1.116296e-09, 
    1.117696e-09, 1.114822e-09, 1.103628e-09, 1.106918e-09, 1.097107e-09, 
    1.091207e-09, 1.087288e-09, 1.084508e-09, 1.084901e-09, 1.08565e-09, 
    1.089501e-09, 1.093122e-09, 1.095881e-09, 1.097727e-09, 1.099546e-09, 
    1.105051e-09, 1.107964e-09, 1.114488e-09, 1.11331e-09, 1.115305e-09, 
    1.11721e-09, 1.120409e-09, 1.119883e-09, 1.121292e-09, 1.115252e-09, 
    1.119266e-09, 1.11264e-09, 1.114452e-09, 1.100041e-09, 1.094549e-09, 
    1.092216e-09, 1.090173e-09, 1.085203e-09, 1.088635e-09, 1.087282e-09, 
    1.090501e-09, 1.092546e-09, 1.091535e-09, 1.097778e-09, 1.09535e-09, 
    1.108137e-09, 1.102629e-09, 1.116988e-09, 1.113552e-09, 1.117812e-09, 
    1.115638e-09, 1.119362e-09, 1.11601e-09, 1.121817e-09, 1.123081e-09, 
    1.122217e-09, 1.125536e-09, 1.115825e-09, 1.119554e-09, 1.091506e-09, 
    1.091671e-09, 1.09244e-09, 1.089061e-09, 1.088855e-09, 1.085758e-09, 
    1.088513e-09, 1.089687e-09, 1.092665e-09, 1.094426e-09, 1.096101e-09, 
    1.099782e-09, 1.103894e-09, 1.109644e-09, 1.113775e-09, 1.116544e-09, 
    1.114846e-09, 1.116345e-09, 1.114669e-09, 1.113884e-09, 1.122607e-09, 
    1.117709e-09, 1.125058e-09, 1.124651e-09, 1.121325e-09, 1.124697e-09, 
    1.091787e-09, 1.090838e-09, 1.087542e-09, 1.090121e-09, 1.085421e-09, 
    1.088052e-09, 1.089565e-09, 1.095401e-09, 1.096683e-09, 1.097873e-09, 
    1.100221e-09, 1.103235e-09, 1.108522e-09, 1.113122e-09, 1.117321e-09, 
    1.117013e-09, 1.117122e-09, 1.11806e-09, 1.115736e-09, 1.118441e-09, 
    1.118895e-09, 1.117708e-09, 1.124597e-09, 1.122629e-09, 1.124643e-09, 
    1.123361e-09, 1.091146e-09, 1.092744e-09, 1.09188e-09, 1.093504e-09, 
    1.09236e-09, 1.097445e-09, 1.09897e-09, 1.106103e-09, 1.103175e-09, 
    1.107835e-09, 1.103649e-09, 1.104391e-09, 1.107987e-09, 1.103875e-09, 
    1.112868e-09, 1.106771e-09, 1.118096e-09, 1.112008e-09, 1.118478e-09, 
    1.117303e-09, 1.119248e-09, 1.12099e-09, 1.123182e-09, 1.127226e-09, 
    1.12629e-09, 1.129672e-09, 1.095125e-09, 1.097197e-09, 1.097015e-09, 
    1.099183e-09, 1.100787e-09, 1.104262e-09, 1.109837e-09, 1.10774e-09, 
    1.111589e-09, 1.112361e-09, 1.106515e-09, 1.110104e-09, 1.098584e-09, 
    1.100445e-09, 1.099337e-09, 1.095289e-09, 1.108224e-09, 1.101585e-09, 
    1.113843e-09, 1.110247e-09, 1.120742e-09, 1.115523e-09, 1.125774e-09, 
    1.130157e-09, 1.134281e-09, 1.139102e-09, 1.098328e-09, 1.09692e-09, 
    1.099441e-09, 1.102929e-09, 1.106164e-09, 1.110466e-09, 1.110906e-09, 
    1.111712e-09, 1.1138e-09, 1.115555e-09, 1.111967e-09, 1.115995e-09, 
    1.100877e-09, 1.1088e-09, 1.096388e-09, 1.100125e-09, 1.102723e-09, 
    1.101583e-09, 1.107501e-09, 1.108895e-09, 1.114563e-09, 1.111633e-09, 
    1.129075e-09, 1.121358e-09, 1.142772e-09, 1.136788e-09, 1.096428e-09, 
    1.098323e-09, 1.104918e-09, 1.10178e-09, 1.110753e-09, 1.112962e-09, 
    1.114758e-09, 1.117053e-09, 1.117301e-09, 1.118661e-09, 1.116432e-09, 
    1.118573e-09, 1.110475e-09, 1.114094e-09, 1.104164e-09, 1.106581e-09, 
    1.105469e-09, 1.104249e-09, 1.108013e-09, 1.112024e-09, 1.112109e-09, 
    1.113395e-09, 1.117019e-09, 1.11079e-09, 1.130072e-09, 1.118164e-09, 
    1.100389e-09, 1.104039e-09, 1.10456e-09, 1.103147e-09, 1.112741e-09, 
    1.109265e-09, 1.118628e-09, 1.116097e-09, 1.120243e-09, 1.118183e-09, 
    1.11788e-09, 1.115234e-09, 1.113586e-09, 1.109424e-09, 1.106037e-09, 
    1.103352e-09, 1.103976e-09, 1.106926e-09, 1.112269e-09, 1.117323e-09, 
    1.116216e-09, 1.119928e-09, 1.110103e-09, 1.114223e-09, 1.112631e-09, 
    1.116783e-09, 1.107685e-09, 1.115433e-09, 1.105704e-09, 1.106557e-09, 
    1.109196e-09, 1.114502e-09, 1.115676e-09, 1.11693e-09, 1.116156e-09, 
    1.112405e-09, 1.11179e-09, 1.109131e-09, 1.108397e-09, 1.106372e-09, 
    1.104694e-09, 1.106227e-09, 1.107836e-09, 1.112406e-09, 1.116525e-09, 
    1.121015e-09, 1.122114e-09, 1.127361e-09, 1.12309e-09, 1.130138e-09, 
    1.124146e-09, 1.134518e-09, 1.115881e-09, 1.12397e-09, 1.109316e-09, 
    1.110894e-09, 1.11375e-09, 1.120299e-09, 1.116763e-09, 1.120898e-09, 
    1.111766e-09, 1.107028e-09, 1.105802e-09, 1.103515e-09, 1.105854e-09, 
    1.105664e-09, 1.107903e-09, 1.107183e-09, 1.112558e-09, 1.109671e-09, 
    1.117872e-09, 1.120865e-09, 1.129317e-09, 1.134499e-09, 1.139773e-09, 
    1.142101e-09, 1.14281e-09, 1.143106e-09 ;

 SOIL2C_TO_SOIL3C =
  7.75817e-11, 7.79231e-11, 7.785673e-11, 7.813209e-11, 7.797934e-11, 
    7.815965e-11, 7.765092e-11, 7.793666e-11, 7.775425e-11, 7.761244e-11, 
    7.866648e-11, 7.814437e-11, 7.920876e-11, 7.887579e-11, 7.97122e-11, 
    7.915694e-11, 7.982415e-11, 7.969617e-11, 8.008135e-11, 7.9971e-11, 
    8.04637e-11, 8.013228e-11, 8.071908e-11, 8.038455e-11, 8.043689e-11, 
    8.012135e-11, 7.824943e-11, 7.860148e-11, 7.822858e-11, 7.827878e-11, 
    7.825626e-11, 7.79825e-11, 7.784455e-11, 7.755561e-11, 7.760807e-11, 
    7.782028e-11, 7.830135e-11, 7.813804e-11, 7.85496e-11, 7.854031e-11, 
    7.89985e-11, 7.879191e-11, 7.9562e-11, 7.934313e-11, 7.997561e-11, 
    7.981655e-11, 7.996814e-11, 7.992217e-11, 7.996874e-11, 7.973546e-11, 
    7.983541e-11, 7.963013e-11, 7.88306e-11, 7.906558e-11, 7.836476e-11, 
    7.794337e-11, 7.766345e-11, 7.746483e-11, 7.749291e-11, 7.754644e-11, 
    7.782152e-11, 7.808014e-11, 7.827723e-11, 7.840907e-11, 7.853897e-11, 
    7.893219e-11, 7.91403e-11, 7.960627e-11, 7.952217e-11, 7.966464e-11, 
    7.980073e-11, 8.002923e-11, 7.999161e-11, 8.009229e-11, 7.966087e-11, 
    7.994759e-11, 7.947427e-11, 7.960373e-11, 7.857432e-11, 7.81821e-11, 
    7.801541e-11, 7.786949e-11, 7.751449e-11, 7.775965e-11, 7.766301e-11, 
    7.789291e-11, 7.803901e-11, 7.796675e-11, 7.841268e-11, 7.823932e-11, 
    7.915263e-11, 7.875924e-11, 7.978485e-11, 7.953943e-11, 7.984368e-11, 
    7.968842e-11, 7.995445e-11, 7.971503e-11, 8.012975e-11, 8.022006e-11, 
    8.015835e-11, 8.03954e-11, 7.970176e-11, 7.996814e-11, 7.796473e-11, 
    7.797651e-11, 7.803141e-11, 7.779009e-11, 7.777533e-11, 7.755417e-11, 
    7.775096e-11, 7.783475e-11, 7.804747e-11, 7.81733e-11, 7.829291e-11, 
    7.85559e-11, 7.88496e-11, 7.926029e-11, 7.955533e-11, 7.975311e-11, 
    7.963184e-11, 7.973891e-11, 7.961921e-11, 7.956312e-11, 8.018622e-11, 
    7.983635e-11, 8.03613e-11, 8.033225e-11, 8.009468e-11, 8.033552e-11, 
    7.798479e-11, 7.791697e-11, 7.768153e-11, 7.786579e-11, 7.753009e-11, 
    7.7718e-11, 7.782605e-11, 7.824295e-11, 7.833453e-11, 7.841947e-11, 
    7.858721e-11, 7.880249e-11, 7.918013e-11, 7.95087e-11, 7.980864e-11, 
    7.978666e-11, 7.97944e-11, 7.986141e-11, 7.969543e-11, 7.988866e-11, 
    7.992109e-11, 7.98363e-11, 8.032836e-11, 8.018778e-11, 8.033163e-11, 
    8.02401e-11, 7.793902e-11, 7.805312e-11, 7.799146e-11, 7.810741e-11, 
    7.802572e-11, 7.838894e-11, 7.849783e-11, 7.900737e-11, 7.879825e-11, 
    7.913106e-11, 7.883205e-11, 7.888504e-11, 7.914193e-11, 7.884821e-11, 
    7.949059e-11, 7.905509e-11, 7.986402e-11, 7.942914e-11, 7.989127e-11, 
    7.980734e-11, 7.994629e-11, 8.007073e-11, 8.022729e-11, 8.051616e-11, 
    8.044927e-11, 8.069084e-11, 7.822323e-11, 7.837123e-11, 7.835819e-11, 
    7.851307e-11, 7.862761e-11, 7.887587e-11, 7.927405e-11, 7.912431e-11, 
    7.939919e-11, 7.945437e-11, 7.903676e-11, 7.929318e-11, 7.847027e-11, 
    7.860324e-11, 7.852406e-11, 7.82349e-11, 7.915883e-11, 7.868467e-11, 
    7.956021e-11, 7.930336e-11, 8.005299e-11, 7.968019e-11, 8.041245e-11, 
    8.07255e-11, 8.102009e-11, 8.13644e-11, 7.845199e-11, 7.835143e-11, 
    7.853149e-11, 7.878061e-11, 7.901174e-11, 7.931902e-11, 7.935046e-11, 
    7.940803e-11, 7.955714e-11, 7.968251e-11, 7.942624e-11, 7.971394e-11, 
    7.863408e-11, 7.919998e-11, 7.831342e-11, 7.858039e-11, 7.876592e-11, 
    7.868453e-11, 7.91072e-11, 7.920681e-11, 7.961163e-11, 7.940237e-11, 
    8.064824e-11, 8.009703e-11, 8.162654e-11, 8.119911e-11, 7.83163e-11, 
    7.845164e-11, 7.892271e-11, 7.869858e-11, 7.933953e-11, 7.94973e-11, 
    7.962556e-11, 7.978952e-11, 7.980721e-11, 7.990435e-11, 7.974517e-11, 
    7.989806e-11, 7.931968e-11, 7.957814e-11, 7.886886e-11, 7.90415e-11, 
    7.896207e-11, 7.887496e-11, 7.914382e-11, 7.943027e-11, 7.943638e-11, 
    7.952823e-11, 7.978709e-11, 7.934213e-11, 8.07194e-11, 7.986885e-11, 
    7.859923e-11, 7.885995e-11, 7.889717e-11, 7.879618e-11, 7.948149e-11, 
    7.923318e-11, 7.990198e-11, 7.972122e-11, 8.001739e-11, 7.987022e-11, 
    7.984857e-11, 7.965955e-11, 7.954187e-11, 7.924457e-11, 7.900266e-11, 
    7.881083e-11, 7.885543e-11, 7.906616e-11, 7.94478e-11, 7.980882e-11, 
    7.972974e-11, 7.999488e-11, 7.929306e-11, 7.958735e-11, 7.947362e-11, 
    7.977018e-11, 7.912034e-11, 7.967375e-11, 7.897888e-11, 7.90398e-11, 
    7.922825e-11, 7.960732e-11, 7.969117e-11, 7.978072e-11, 7.972546e-11, 
    7.945748e-11, 7.941357e-11, 7.922367e-11, 7.917124e-11, 7.902654e-11, 
    7.890674e-11, 7.90162e-11, 7.913115e-11, 7.945759e-11, 7.975177e-11, 
    8.007251e-11, 8.0151e-11, 8.052577e-11, 8.022071e-11, 8.072414e-11, 
    8.029614e-11, 8.103701e-11, 7.97058e-11, 8.028354e-11, 7.923683e-11, 
    7.934959e-11, 7.955355e-11, 8.002134e-11, 7.976879e-11, 8.006415e-11, 
    7.941185e-11, 7.907343e-11, 7.898586e-11, 7.882249e-11, 7.898959e-11, 
    7.8976e-11, 7.91359e-11, 7.908452e-11, 7.946842e-11, 7.926221e-11, 
    7.984803e-11, 8.006181e-11, 8.066553e-11, 8.103563e-11, 8.141236e-11, 
    8.157867e-11, 8.16293e-11, 8.165046e-11 ;

 SOIL2C_vr =
  20.00646, 20.00648, 20.00648, 20.00649, 20.00648, 20.00649, 20.00646, 
    20.00648, 20.00647, 20.00646, 20.00652, 20.00649, 20.00654, 20.00653, 
    20.00657, 20.00654, 20.00657, 20.00657, 20.00658, 20.00658, 20.0066, 
    20.00659, 20.00661, 20.0066, 20.0066, 20.00659, 20.00649, 20.00651, 
    20.00649, 20.0065, 20.00649, 20.00648, 20.00647, 20.00646, 20.00646, 
    20.00647, 20.0065, 20.00649, 20.00651, 20.00651, 20.00653, 20.00652, 
    20.00656, 20.00655, 20.00658, 20.00657, 20.00658, 20.00658, 20.00658, 
    20.00657, 20.00657, 20.00656, 20.00652, 20.00653, 20.0065, 20.00648, 
    20.00647, 20.00646, 20.00646, 20.00646, 20.00647, 20.00649, 20.0065, 
    20.0065, 20.00651, 20.00653, 20.00654, 20.00656, 20.00656, 20.00656, 
    20.00657, 20.00658, 20.00658, 20.00658, 20.00656, 20.00658, 20.00656, 
    20.00656, 20.00651, 20.00649, 20.00648, 20.00648, 20.00646, 20.00647, 
    20.00647, 20.00648, 20.00648, 20.00648, 20.0065, 20.00649, 20.00654, 
    20.00652, 20.00657, 20.00656, 20.00657, 20.00657, 20.00658, 20.00657, 
    20.00659, 20.00659, 20.00659, 20.0066, 20.00657, 20.00658, 20.00648, 
    20.00648, 20.00648, 20.00647, 20.00647, 20.00646, 20.00647, 20.00647, 
    20.00648, 20.00649, 20.0065, 20.00651, 20.00652, 20.00654, 20.00656, 
    20.00657, 20.00656, 20.00657, 20.00656, 20.00656, 20.00659, 20.00657, 
    20.0066, 20.0066, 20.00658, 20.0066, 20.00648, 20.00648, 20.00647, 
    20.00648, 20.00646, 20.00647, 20.00647, 20.00649, 20.0065, 20.0065, 
    20.00651, 20.00652, 20.00654, 20.00656, 20.00657, 20.00657, 20.00657, 
    20.00657, 20.00657, 20.00657, 20.00658, 20.00657, 20.0066, 20.00659, 
    20.0066, 20.00659, 20.00648, 20.00648, 20.00648, 20.00649, 20.00648, 
    20.0065, 20.00651, 20.00653, 20.00652, 20.00654, 20.00652, 20.00653, 
    20.00654, 20.00652, 20.00656, 20.00653, 20.00657, 20.00655, 20.00657, 
    20.00657, 20.00658, 20.00658, 20.00659, 20.00661, 20.0066, 20.00661, 
    20.00649, 20.0065, 20.0065, 20.00651, 20.00651, 20.00653, 20.00654, 
    20.00654, 20.00655, 20.00655, 20.00653, 20.00655, 20.00651, 20.00651, 
    20.00651, 20.00649, 20.00654, 20.00652, 20.00656, 20.00655, 20.00658, 
    20.00657, 20.0066, 20.00662, 20.00663, 20.00665, 20.0065, 20.0065, 
    20.00651, 20.00652, 20.00653, 20.00655, 20.00655, 20.00655, 20.00656, 
    20.00657, 20.00655, 20.00657, 20.00651, 20.00654, 20.0065, 20.00651, 
    20.00652, 20.00652, 20.00654, 20.00654, 20.00656, 20.00655, 20.00661, 
    20.00659, 20.00666, 20.00664, 20.0065, 20.0065, 20.00653, 20.00652, 
    20.00655, 20.00656, 20.00656, 20.00657, 20.00657, 20.00658, 20.00657, 
    20.00657, 20.00655, 20.00656, 20.00653, 20.00653, 20.00653, 20.00653, 
    20.00654, 20.00655, 20.00655, 20.00656, 20.00657, 20.00655, 20.00662, 
    20.00657, 20.00651, 20.00653, 20.00653, 20.00652, 20.00656, 20.00654, 
    20.00658, 20.00657, 20.00658, 20.00657, 20.00657, 20.00656, 20.00656, 
    20.00654, 20.00653, 20.00652, 20.00653, 20.00653, 20.00655, 20.00657, 
    20.00657, 20.00658, 20.00655, 20.00656, 20.00655, 20.00657, 20.00654, 
    20.00657, 20.00653, 20.00653, 20.00654, 20.00656, 20.00657, 20.00657, 
    20.00657, 20.00655, 20.00655, 20.00654, 20.00654, 20.00653, 20.00653, 
    20.00653, 20.00654, 20.00655, 20.00657, 20.00658, 20.00659, 20.00661, 
    20.00659, 20.00662, 20.0066, 20.00663, 20.00657, 20.00659, 20.00654, 
    20.00655, 20.00656, 20.00658, 20.00657, 20.00658, 20.00655, 20.00653, 
    20.00653, 20.00652, 20.00653, 20.00653, 20.00654, 20.00653, 20.00655, 
    20.00654, 20.00657, 20.00658, 20.00661, 20.00663, 20.00665, 20.00666, 
    20.00666, 20.00666,
  20.00607, 20.00609, 20.00609, 20.00611, 20.0061, 20.00611, 20.00607, 
    20.00609, 20.00608, 20.00607, 20.00614, 20.00611, 20.00618, 20.00616, 
    20.00621, 20.00617, 20.00622, 20.00621, 20.00624, 20.00623, 20.00626, 
    20.00624, 20.00628, 20.00626, 20.00626, 20.00624, 20.00611, 20.00614, 
    20.00611, 20.00612, 20.00611, 20.0061, 20.00609, 20.00607, 20.00607, 
    20.00609, 20.00612, 20.00611, 20.00613, 20.00613, 20.00616, 20.00615, 
    20.0062, 20.00619, 20.00623, 20.00622, 20.00623, 20.00623, 20.00623, 
    20.00621, 20.00622, 20.00621, 20.00615, 20.00617, 20.00612, 20.00609, 
    20.00607, 20.00606, 20.00606, 20.00607, 20.00609, 20.0061, 20.00612, 
    20.00612, 20.00613, 20.00616, 20.00617, 20.0062, 20.0062, 20.00621, 
    20.00622, 20.00623, 20.00623, 20.00624, 20.00621, 20.00623, 20.0062, 
    20.0062, 20.00614, 20.00611, 20.0061, 20.00609, 20.00607, 20.00608, 
    20.00607, 20.00609, 20.0061, 20.0061, 20.00612, 20.00611, 20.00617, 
    20.00615, 20.00622, 20.0062, 20.00622, 20.00621, 20.00623, 20.00621, 
    20.00624, 20.00624, 20.00624, 20.00626, 20.00621, 20.00623, 20.0061, 
    20.0061, 20.0061, 20.00608, 20.00608, 20.00607, 20.00608, 20.00609, 
    20.0061, 20.00611, 20.00612, 20.00613, 20.00615, 20.00618, 20.0062, 
    20.00621, 20.00621, 20.00621, 20.0062, 20.0062, 20.00624, 20.00622, 
    20.00625, 20.00625, 20.00624, 20.00625, 20.0061, 20.00609, 20.00608, 
    20.00609, 20.00607, 20.00608, 20.00609, 20.00611, 20.00612, 20.00612, 
    20.00614, 20.00615, 20.00618, 20.0062, 20.00622, 20.00622, 20.00622, 
    20.00622, 20.00621, 20.00622, 20.00623, 20.00622, 20.00625, 20.00624, 
    20.00625, 20.00625, 20.00609, 20.0061, 20.0061, 20.00611, 20.0061, 
    20.00612, 20.00613, 20.00616, 20.00615, 20.00617, 20.00615, 20.00616, 
    20.00617, 20.00615, 20.0062, 20.00617, 20.00622, 20.00619, 20.00622, 
    20.00622, 20.00623, 20.00624, 20.00624, 20.00626, 20.00626, 20.00628, 
    20.00611, 20.00612, 20.00612, 20.00613, 20.00614, 20.00616, 20.00618, 
    20.00617, 20.00619, 20.00619, 20.00617, 20.00618, 20.00613, 20.00614, 
    20.00613, 20.00611, 20.00617, 20.00614, 20.0062, 20.00618, 20.00623, 
    20.00621, 20.00626, 20.00628, 20.0063, 20.00632, 20.00613, 20.00612, 
    20.00613, 20.00615, 20.00616, 20.00619, 20.00619, 20.00619, 20.0062, 
    20.00621, 20.00619, 20.00621, 20.00614, 20.00618, 20.00612, 20.00614, 
    20.00615, 20.00614, 20.00617, 20.00618, 20.0062, 20.00619, 20.00627, 
    20.00624, 20.00634, 20.00631, 20.00612, 20.00613, 20.00616, 20.00614, 
    20.00619, 20.0062, 20.0062, 20.00622, 20.00622, 20.00622, 20.00621, 
    20.00622, 20.00619, 20.0062, 20.00616, 20.00617, 20.00616, 20.00616, 
    20.00617, 20.00619, 20.00619, 20.0062, 20.00622, 20.00619, 20.00628, 
    20.00622, 20.00614, 20.00616, 20.00616, 20.00615, 20.0062, 20.00618, 
    20.00622, 20.00621, 20.00623, 20.00622, 20.00622, 20.00621, 20.0062, 
    20.00618, 20.00616, 20.00615, 20.00616, 20.00617, 20.00619, 20.00622, 
    20.00621, 20.00623, 20.00618, 20.0062, 20.0062, 20.00621, 20.00617, 
    20.00621, 20.00616, 20.00617, 20.00618, 20.0062, 20.00621, 20.00622, 
    20.00621, 20.0062, 20.00619, 20.00618, 20.00618, 20.00617, 20.00616, 
    20.00616, 20.00617, 20.0062, 20.00621, 20.00624, 20.00624, 20.00627, 
    20.00624, 20.00628, 20.00625, 20.0063, 20.00621, 20.00625, 20.00618, 
    20.00619, 20.0062, 20.00623, 20.00621, 20.00624, 20.00619, 20.00617, 
    20.00616, 20.00615, 20.00616, 20.00616, 20.00617, 20.00617, 20.0062, 
    20.00618, 20.00622, 20.00623, 20.00627, 20.0063, 20.00632, 20.00633, 
    20.00634, 20.00634,
  20.00552, 20.00554, 20.00554, 20.00556, 20.00555, 20.00556, 20.00552, 
    20.00554, 20.00553, 20.00552, 20.0056, 20.00556, 20.00563, 20.00561, 
    20.00567, 20.00563, 20.00568, 20.00567, 20.0057, 20.00569, 20.00572, 
    20.0057, 20.00574, 20.00572, 20.00572, 20.0057, 20.00557, 20.00559, 
    20.00557, 20.00557, 20.00557, 20.00555, 20.00554, 20.00552, 20.00552, 
    20.00554, 20.00557, 20.00556, 20.00559, 20.00559, 20.00562, 20.00561, 
    20.00566, 20.00564, 20.00569, 20.00568, 20.00569, 20.00569, 20.00569, 
    20.00567, 20.00568, 20.00566, 20.00561, 20.00562, 20.00558, 20.00554, 
    20.00553, 20.00551, 20.00551, 20.00552, 20.00554, 20.00555, 20.00557, 
    20.00558, 20.00559, 20.00562, 20.00563, 20.00566, 20.00566, 20.00567, 
    20.00568, 20.00569, 20.00569, 20.0057, 20.00567, 20.00569, 20.00565, 
    20.00566, 20.00559, 20.00556, 20.00555, 20.00554, 20.00551, 20.00553, 
    20.00553, 20.00554, 20.00555, 20.00555, 20.00558, 20.00557, 20.00563, 
    20.0056, 20.00567, 20.00566, 20.00568, 20.00567, 20.00569, 20.00567, 
    20.0057, 20.00571, 20.0057, 20.00572, 20.00567, 20.00569, 20.00555, 
    20.00555, 20.00555, 20.00553, 20.00553, 20.00552, 20.00553, 20.00554, 
    20.00555, 20.00556, 20.00557, 20.00559, 20.00561, 20.00564, 20.00566, 
    20.00567, 20.00566, 20.00567, 20.00566, 20.00566, 20.0057, 20.00568, 
    20.00572, 20.00571, 20.0057, 20.00571, 20.00555, 20.00554, 20.00553, 
    20.00554, 20.00552, 20.00553, 20.00554, 20.00557, 20.00557, 20.00558, 
    20.00559, 20.00561, 20.00563, 20.00566, 20.00568, 20.00568, 20.00568, 
    20.00568, 20.00567, 20.00568, 20.00569, 20.00568, 20.00571, 20.0057, 
    20.00571, 20.00571, 20.00554, 20.00555, 20.00555, 20.00556, 20.00555, 
    20.00558, 20.00558, 20.00562, 20.00561, 20.00563, 20.00561, 20.00561, 
    20.00563, 20.00561, 20.00566, 20.00562, 20.00568, 20.00565, 20.00568, 
    20.00568, 20.00569, 20.0057, 20.00571, 20.00573, 20.00572, 20.00574, 
    20.00557, 20.00558, 20.00558, 20.00558, 20.00559, 20.00561, 20.00564, 
    20.00563, 20.00565, 20.00565, 20.00562, 20.00564, 20.00558, 20.00559, 
    20.00559, 20.00557, 20.00563, 20.0056, 20.00566, 20.00564, 20.00569, 
    20.00567, 20.00572, 20.00574, 20.00576, 20.00579, 20.00558, 20.00557, 
    20.00559, 20.0056, 20.00562, 20.00564, 20.00564, 20.00565, 20.00566, 
    20.00567, 20.00565, 20.00567, 20.00559, 20.00563, 20.00557, 20.00559, 
    20.0056, 20.0056, 20.00563, 20.00563, 20.00566, 20.00565, 20.00574, 
    20.0057, 20.00581, 20.00578, 20.00557, 20.00558, 20.00562, 20.0056, 
    20.00564, 20.00566, 20.00566, 20.00568, 20.00568, 20.00568, 20.00567, 
    20.00568, 20.00564, 20.00566, 20.00561, 20.00562, 20.00562, 20.00561, 
    20.00563, 20.00565, 20.00565, 20.00566, 20.00568, 20.00564, 20.00574, 
    20.00568, 20.00559, 20.00561, 20.00561, 20.00561, 20.00565, 20.00564, 
    20.00568, 20.00567, 20.00569, 20.00568, 20.00568, 20.00567, 20.00566, 
    20.00564, 20.00562, 20.00561, 20.00561, 20.00562, 20.00565, 20.00568, 
    20.00567, 20.00569, 20.00564, 20.00566, 20.00565, 20.00567, 20.00563, 
    20.00567, 20.00562, 20.00562, 20.00564, 20.00566, 20.00567, 20.00567, 
    20.00567, 20.00565, 20.00565, 20.00564, 20.00563, 20.00562, 20.00561, 
    20.00562, 20.00563, 20.00565, 20.00567, 20.0057, 20.0057, 20.00573, 
    20.00571, 20.00574, 20.00571, 20.00576, 20.00567, 20.00571, 20.00564, 
    20.00564, 20.00566, 20.00569, 20.00567, 20.0057, 20.00565, 20.00562, 
    20.00562, 20.00561, 20.00562, 20.00562, 20.00563, 20.00563, 20.00565, 
    20.00564, 20.00568, 20.0057, 20.00574, 20.00576, 20.00579, 20.0058, 
    20.00581, 20.00581,
  20.00508, 20.0051, 20.0051, 20.00512, 20.00511, 20.00512, 20.00508, 
    20.00511, 20.00509, 20.00508, 20.00516, 20.00512, 20.00519, 20.00517, 
    20.00523, 20.00519, 20.00524, 20.00523, 20.00525, 20.00525, 20.00528, 
    20.00526, 20.0053, 20.00528, 20.00528, 20.00526, 20.00513, 20.00515, 
    20.00513, 20.00513, 20.00513, 20.00511, 20.0051, 20.00508, 20.00508, 
    20.0051, 20.00513, 20.00512, 20.00515, 20.00515, 20.00518, 20.00517, 
    20.00522, 20.0052, 20.00525, 20.00524, 20.00525, 20.00525, 20.00525, 
    20.00523, 20.00524, 20.00522, 20.00517, 20.00518, 20.00513, 20.00511, 
    20.00508, 20.00507, 20.00507, 20.00508, 20.0051, 20.00512, 20.00513, 
    20.00514, 20.00515, 20.00517, 20.00519, 20.00522, 20.00522, 20.00523, 
    20.00524, 20.00525, 20.00525, 20.00526, 20.00523, 20.00525, 20.00521, 
    20.00522, 20.00515, 20.00512, 20.00511, 20.0051, 20.00508, 20.00509, 
    20.00508, 20.0051, 20.00511, 20.00511, 20.00514, 20.00513, 20.00519, 
    20.00516, 20.00524, 20.00522, 20.00524, 20.00523, 20.00525, 20.00523, 
    20.00526, 20.00527, 20.00526, 20.00528, 20.00523, 20.00525, 20.00511, 
    20.00511, 20.00511, 20.00509, 20.00509, 20.00508, 20.00509, 20.0051, 
    20.00511, 20.00512, 20.00513, 20.00515, 20.00517, 20.0052, 20.00522, 
    20.00523, 20.00522, 20.00523, 20.00522, 20.00522, 20.00526, 20.00524, 
    20.00528, 20.00527, 20.00526, 20.00527, 20.00511, 20.0051, 20.00509, 
    20.0051, 20.00508, 20.00509, 20.0051, 20.00513, 20.00513, 20.00514, 
    20.00515, 20.00517, 20.00519, 20.00521, 20.00524, 20.00524, 20.00524, 
    20.00524, 20.00523, 20.00524, 20.00525, 20.00524, 20.00527, 20.00526, 
    20.00527, 20.00527, 20.00511, 20.00511, 20.00511, 20.00512, 20.00511, 
    20.00514, 20.00514, 20.00518, 20.00517, 20.00519, 20.00517, 20.00517, 
    20.00519, 20.00517, 20.00521, 20.00518, 20.00524, 20.00521, 20.00524, 
    20.00524, 20.00525, 20.00525, 20.00527, 20.00529, 20.00528, 20.0053, 
    20.00513, 20.00514, 20.00513, 20.00515, 20.00515, 20.00517, 20.0052, 
    20.00519, 20.00521, 20.00521, 20.00518, 20.0052, 20.00514, 20.00515, 
    20.00515, 20.00513, 20.00519, 20.00516, 20.00522, 20.0052, 20.00525, 
    20.00523, 20.00528, 20.0053, 20.00532, 20.00535, 20.00514, 20.00513, 
    20.00515, 20.00517, 20.00518, 20.0052, 20.00521, 20.00521, 20.00522, 
    20.00523, 20.00521, 20.00523, 20.00515, 20.00519, 20.00513, 20.00515, 
    20.00516, 20.00516, 20.00519, 20.00519, 20.00522, 20.00521, 20.00529, 
    20.00526, 20.00536, 20.00533, 20.00513, 20.00514, 20.00517, 20.00516, 
    20.0052, 20.00521, 20.00522, 20.00524, 20.00524, 20.00524, 20.00523, 
    20.00524, 20.0052, 20.00522, 20.00517, 20.00518, 20.00518, 20.00517, 
    20.00519, 20.00521, 20.00521, 20.00522, 20.00524, 20.0052, 20.0053, 
    20.00524, 20.00515, 20.00517, 20.00517, 20.00517, 20.00521, 20.0052, 
    20.00524, 20.00523, 20.00525, 20.00524, 20.00524, 20.00523, 20.00522, 
    20.0052, 20.00518, 20.00517, 20.00517, 20.00518, 20.00521, 20.00524, 
    20.00523, 20.00525, 20.0052, 20.00522, 20.00521, 20.00523, 20.00519, 
    20.00523, 20.00518, 20.00518, 20.0052, 20.00522, 20.00523, 20.00523, 
    20.00523, 20.00521, 20.00521, 20.0052, 20.00519, 20.00518, 20.00517, 
    20.00518, 20.00519, 20.00521, 20.00523, 20.00525, 20.00526, 20.00529, 
    20.00527, 20.0053, 20.00527, 20.00532, 20.00523, 20.00527, 20.0052, 
    20.00521, 20.00522, 20.00525, 20.00523, 20.00525, 20.00521, 20.00518, 
    20.00518, 20.00517, 20.00518, 20.00518, 20.00519, 20.00519, 20.00521, 
    20.0052, 20.00524, 20.00525, 20.0053, 20.00532, 20.00535, 20.00536, 
    20.00536, 20.00537,
  20.00437, 20.00439, 20.00439, 20.0044, 20.00439, 20.00441, 20.00438, 
    20.00439, 20.00438, 20.00437, 20.00444, 20.0044, 20.00447, 20.00445, 
    20.0045, 20.00447, 20.00451, 20.0045, 20.00452, 20.00451, 20.00454, 
    20.00452, 20.00456, 20.00454, 20.00454, 20.00452, 20.00441, 20.00443, 
    20.00441, 20.00441, 20.00441, 20.00439, 20.00439, 20.00437, 20.00437, 
    20.00438, 20.00441, 20.0044, 20.00443, 20.00443, 20.00446, 20.00444, 
    20.00449, 20.00448, 20.00451, 20.00451, 20.00451, 20.00451, 20.00451, 
    20.0045, 20.00451, 20.00449, 20.00445, 20.00446, 20.00442, 20.00439, 
    20.00438, 20.00436, 20.00437, 20.00437, 20.00438, 20.0044, 20.00441, 
    20.00442, 20.00443, 20.00445, 20.00446, 20.00449, 20.00449, 20.0045, 
    20.0045, 20.00452, 20.00451, 20.00452, 20.0045, 20.00451, 20.00448, 
    20.00449, 20.00443, 20.00441, 20.0044, 20.00439, 20.00437, 20.00438, 
    20.00438, 20.00439, 20.0044, 20.00439, 20.00442, 20.00441, 20.00447, 
    20.00444, 20.0045, 20.00449, 20.00451, 20.0045, 20.00451, 20.0045, 
    20.00452, 20.00453, 20.00452, 20.00454, 20.0045, 20.00451, 20.00439, 
    20.00439, 20.0044, 20.00438, 20.00438, 20.00437, 20.00438, 20.00439, 
    20.0044, 20.00441, 20.00441, 20.00443, 20.00445, 20.00447, 20.00449, 
    20.0045, 20.00449, 20.0045, 20.00449, 20.00449, 20.00453, 20.00451, 
    20.00454, 20.00454, 20.00452, 20.00454, 20.00439, 20.00439, 20.00438, 
    20.00439, 20.00437, 20.00438, 20.00438, 20.00441, 20.00442, 20.00442, 
    20.00443, 20.00444, 20.00447, 20.00449, 20.0045, 20.0045, 20.0045, 
    20.00451, 20.0045, 20.00451, 20.00451, 20.00451, 20.00454, 20.00453, 
    20.00454, 20.00453, 20.00439, 20.0044, 20.00439, 20.0044, 20.0044, 
    20.00442, 20.00443, 20.00446, 20.00444, 20.00446, 20.00445, 20.00445, 
    20.00446, 20.00445, 20.00448, 20.00446, 20.00451, 20.00448, 20.00451, 
    20.0045, 20.00451, 20.00452, 20.00453, 20.00455, 20.00454, 20.00456, 
    20.00441, 20.00442, 20.00442, 20.00443, 20.00443, 20.00445, 20.00447, 
    20.00446, 20.00448, 20.00448, 20.00446, 20.00447, 20.00442, 20.00443, 
    20.00443, 20.00441, 20.00447, 20.00444, 20.00449, 20.00447, 20.00452, 
    20.0045, 20.00454, 20.00456, 20.00458, 20.0046, 20.00442, 20.00442, 
    20.00443, 20.00444, 20.00446, 20.00447, 20.00448, 20.00448, 20.00449, 
    20.0045, 20.00448, 20.0045, 20.00443, 20.00447, 20.00442, 20.00443, 
    20.00444, 20.00444, 20.00446, 20.00447, 20.00449, 20.00448, 20.00455, 
    20.00452, 20.00461, 20.00459, 20.00442, 20.00442, 20.00445, 20.00444, 
    20.00448, 20.00449, 20.00449, 20.0045, 20.0045, 20.00451, 20.0045, 
    20.00451, 20.00447, 20.00449, 20.00445, 20.00446, 20.00445, 20.00445, 
    20.00446, 20.00448, 20.00448, 20.00449, 20.0045, 20.00448, 20.00456, 
    20.00451, 20.00443, 20.00445, 20.00445, 20.00444, 20.00448, 20.00447, 
    20.00451, 20.0045, 20.00452, 20.00451, 20.00451, 20.0045, 20.00449, 
    20.00447, 20.00446, 20.00444, 20.00445, 20.00446, 20.00448, 20.0045, 
    20.0045, 20.00451, 20.00447, 20.00449, 20.00448, 20.0045, 20.00446, 
    20.0045, 20.00445, 20.00446, 20.00447, 20.00449, 20.0045, 20.0045, 
    20.0045, 20.00448, 20.00448, 20.00447, 20.00447, 20.00446, 20.00445, 
    20.00446, 20.00446, 20.00448, 20.0045, 20.00452, 20.00452, 20.00455, 
    20.00453, 20.00456, 20.00453, 20.00458, 20.0045, 20.00453, 20.00447, 
    20.00448, 20.00449, 20.00452, 20.0045, 20.00452, 20.00448, 20.00446, 
    20.00446, 20.00444, 20.00446, 20.00445, 20.00446, 20.00446, 20.00448, 
    20.00447, 20.00451, 20.00452, 20.00455, 20.00458, 20.0046, 20.00461, 
    20.00461, 20.00461,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N =
  0.5258222, 0.5258228, 0.5258227, 0.5258232, 0.5258229, 0.5258232, 
    0.5258223, 0.5258228, 0.5258225, 0.5258223, 0.5258241, 0.5258232, 
    0.525825, 0.5258244, 0.5258258, 0.5258249, 0.525826, 0.5258258, 
    0.5258265, 0.5258263, 0.5258271, 0.5258265, 0.5258275, 0.5258269, 
    0.5258271, 0.5258265, 0.5258234, 0.525824, 0.5258233, 0.5258234, 
    0.5258234, 0.5258229, 0.5258227, 0.5258222, 0.5258223, 0.5258226, 
    0.5258235, 0.5258232, 0.5258239, 0.5258238, 0.5258246, 0.5258242, 
    0.5258256, 0.5258252, 0.5258263, 0.525826, 0.5258263, 0.5258262, 
    0.5258263, 0.5258259, 0.525826, 0.5258257, 0.5258243, 0.5258247, 
    0.5258235, 0.5258228, 0.5258223, 0.525822, 0.5258221, 0.5258222, 
    0.5258226, 0.5258231, 0.5258234, 0.5258237, 0.5258238, 0.5258245, 
    0.5258248, 0.5258256, 0.5258255, 0.5258257, 0.525826, 0.5258263, 
    0.5258263, 0.5258265, 0.5258257, 0.5258262, 0.5258254, 0.5258256, 
    0.5258239, 0.5258232, 0.5258229, 0.5258227, 0.5258221, 0.5258225, 
    0.5258223, 0.5258228, 0.525823, 0.5258229, 0.5258237, 0.5258234, 
    0.5258249, 0.5258242, 0.5258259, 0.5258256, 0.525826, 0.5258258, 
    0.5258262, 0.5258258, 0.5258265, 0.5258267, 0.5258266, 0.525827, 
    0.5258258, 0.5258263, 0.5258229, 0.5258229, 0.525823, 0.5258226, 
    0.5258226, 0.5258222, 0.5258225, 0.5258226, 0.525823, 0.5258232, 
    0.5258234, 0.5258239, 0.5258244, 0.5258251, 0.5258256, 0.5258259, 
    0.5258257, 0.5258259, 0.5258257, 0.5258256, 0.5258266, 0.525826, 
    0.5258269, 0.5258269, 0.5258265, 0.5258269, 0.5258229, 0.5258228, 
    0.5258224, 0.5258227, 0.5258222, 0.5258225, 0.5258226, 0.5258234, 
    0.5258235, 0.5258237, 0.525824, 0.5258243, 0.5258249, 0.5258255, 
    0.525826, 0.525826, 0.525826, 0.5258261, 0.5258258, 0.5258261, 0.5258262, 
    0.525826, 0.5258269, 0.5258266, 0.5258269, 0.5258267, 0.5258228, 
    0.525823, 0.5258229, 0.5258231, 0.525823, 0.5258236, 0.5258238, 
    0.5258246, 0.5258243, 0.5258248, 0.5258244, 0.5258244, 0.5258248, 
    0.5258244, 0.5258254, 0.5258247, 0.5258261, 0.5258253, 0.5258261, 
    0.525826, 0.5258262, 0.5258265, 0.5258267, 0.5258272, 0.5258271, 
    0.5258275, 0.5258233, 0.5258235, 0.5258235, 0.5258238, 0.525824, 
    0.5258244, 0.5258251, 0.5258248, 0.5258253, 0.5258254, 0.5258247, 
    0.5258251, 0.5258237, 0.525824, 0.5258238, 0.5258234, 0.5258249, 
    0.5258241, 0.5258256, 0.5258251, 0.5258264, 0.5258258, 0.525827, 
    0.5258275, 0.525828, 0.5258286, 0.5258237, 0.5258235, 0.5258238, 
    0.5258242, 0.5258247, 0.5258251, 0.5258252, 0.5258253, 0.5258256, 
    0.5258258, 0.5258253, 0.5258258, 0.525824, 0.525825, 0.5258235, 
    0.5258239, 0.5258242, 0.5258241, 0.5258248, 0.525825, 0.5258257, 
    0.5258253, 0.5258274, 0.5258265, 0.5258291, 0.5258283, 0.5258235, 
    0.5258237, 0.5258245, 0.5258241, 0.5258252, 0.5258254, 0.5258257, 
    0.525826, 0.525826, 0.5258262, 0.5258259, 0.5258262, 0.5258251, 
    0.5258256, 0.5258244, 0.5258247, 0.5258245, 0.5258244, 0.5258248, 
    0.5258253, 0.5258254, 0.5258255, 0.525826, 0.5258252, 0.5258275, 
    0.5258261, 0.525824, 0.5258244, 0.5258244, 0.5258243, 0.5258254, 
    0.525825, 0.5258262, 0.5258259, 0.5258263, 0.5258261, 0.525826, 
    0.5258257, 0.5258256, 0.525825, 0.5258246, 0.5258243, 0.5258244, 
    0.5258247, 0.5258254, 0.525826, 0.5258259, 0.5258263, 0.5258251, 
    0.5258256, 0.5258254, 0.5258259, 0.5258248, 0.5258257, 0.5258246, 
    0.5258247, 0.525825, 0.5258256, 0.5258258, 0.5258259, 0.5258259, 
    0.5258254, 0.5258253, 0.525825, 0.5258249, 0.5258247, 0.5258245, 
    0.5258247, 0.5258248, 0.5258254, 0.5258259, 0.5258265, 0.5258266, 
    0.5258272, 0.5258267, 0.5258275, 0.5258268, 0.5258281, 0.5258258, 
    0.5258268, 0.525825, 0.5258252, 0.5258256, 0.5258263, 0.5258259, 
    0.5258264, 0.5258253, 0.5258247, 0.5258246, 0.5258243, 0.5258246, 
    0.5258246, 0.5258248, 0.5258248, 0.5258254, 0.5258251, 0.525826, 
    0.5258264, 0.5258274, 0.5258281, 0.5258287, 0.525829, 0.5258291, 0.5258291 ;

 SOIL2N_TNDNCY_VERT_TRANS =
  -1.798972e-20, -1.798972e-20, -7.709882e-21, 2.569961e-21, -5.139921e-21, 
    -1.541976e-20, -5.139921e-21, 7.709882e-21, 0, -2.569961e-21, 
    -1.28498e-20, -5.139921e-21, 5.139921e-21, 1.28498e-20, 1.28498e-20, 
    -2.312965e-20, -5.139921e-21, -7.709882e-21, -1.027984e-20, 2.569961e-21, 
    -2.569961e-21, -2.569961e-21, 2.055969e-20, -7.709882e-21, 1.003089e-36, 
    -2.569961e-21, 5.139921e-21, 2.569961e-21, -2.569961e-21, -1.541976e-20, 
    -1.541976e-20, -2.569961e-21, 7.709882e-21, -5.139921e-21, -2.569961e-21, 
    7.709882e-21, 2.569961e-21, -1.027984e-20, -2.569961e-21, -5.139921e-21, 
    5.139921e-21, 1.541976e-20, 5.139921e-21, -1.28498e-20, -1.027984e-20, 
    2.569961e-21, -1.027984e-20, -2.569961e-21, 5.139921e-21, -1.798972e-20, 
    -7.709882e-21, -7.709882e-21, -1.027984e-20, 1.28498e-20, -1.541976e-20, 
    2.569961e-20, -5.139921e-21, 5.139921e-21, 2.569961e-21, -5.139921e-21, 
    5.139921e-21, 0, 2.569961e-21, -1.28498e-20, -5.139921e-21, 
    -7.709882e-21, 7.709882e-21, -1.541976e-20, 2.569961e-21, -1.027984e-20, 
    1.798972e-20, 5.139921e-21, -1.541976e-20, 5.139921e-21, -1.003089e-36, 
    -7.709882e-21, 5.139921e-21, 1.027984e-20, 1.003089e-36, 2.569961e-21, 
    1.28498e-20, 5.139921e-21, 2.569961e-21, 0, 1.798972e-20, -5.139921e-21, 
    2.569961e-21, 0, 1.798972e-20, -2.055969e-20, 1.027984e-20, 5.139921e-21, 
    7.709882e-21, 1.003089e-36, -2.312965e-20, -5.139921e-21, -2.312965e-20, 
    -7.709882e-21, 5.139921e-21, 1.541976e-20, -1.28498e-20, 7.709882e-21, 
    5.139921e-21, -2.569961e-21, -1.027984e-20, 2.569961e-21, 0, 
    -1.798972e-20, 1.541976e-20, 5.139921e-21, -7.709882e-21, -2.569961e-21, 
    -1.027984e-20, 1.541976e-20, -7.709882e-21, 1.541976e-20, -5.139921e-21, 
    1.541976e-20, -1.541976e-20, 1.027984e-20, 2.569961e-21, -2.569961e-21, 
    7.709882e-21, -1.541976e-20, -1.003089e-36, -1.003089e-36, -1.003089e-36, 
    1.003089e-36, -5.139921e-21, 1.541976e-20, 2.055969e-20, -2.569961e-21, 
    1.28498e-20, 2.569961e-21, -7.709882e-21, 2.569961e-21, 5.139921e-21, 
    1.003089e-36, -2.569961e-21, -2.569961e-21, 2.569961e-21, -1.003089e-36, 
    1.28498e-20, 7.709882e-21, 5.139921e-21, -5.139921e-21, 2.569961e-21, 
    -2.569961e-21, -2.569961e-21, -1.28498e-20, 1.28498e-20, 7.709882e-21, 
    2.312965e-20, 1.798972e-20, 7.709882e-21, -1.798972e-20, -1.003089e-36, 
    1.541976e-20, -2.569961e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    1.003089e-36, 0, -1.027984e-20, -1.798972e-20, -2.569961e-21, 
    -2.569961e-21, 0, -2.569961e-21, -2.569961e-21, 1.027984e-20, 0, 
    3.083953e-20, -2.569961e-21, 2.569961e-21, 7.709882e-21, 1.798972e-20, 
    -2.569961e-21, -1.003089e-36, 7.709882e-21, -1.541976e-20, 2.569961e-21, 
    1.003089e-36, -7.709882e-21, -1.798972e-20, 5.139921e-21, 0, 
    5.139921e-21, 1.027984e-20, 5.139921e-21, 1.28498e-20, -1.027984e-20, 
    1.28498e-20, -7.709882e-21, 7.709882e-21, 2.055969e-20, -1.027984e-20, 
    -5.139921e-21, -1.003089e-36, -5.139921e-21, -5.139921e-21, 2.569961e-21, 
    -1.003089e-36, -1.28498e-20, 1.003089e-36, 1.027984e-20, -1.027984e-20, 
    -5.139921e-21, 5.139921e-21, 1.28498e-20, -1.027984e-20, 1.28498e-20, 
    -1.28498e-20, -7.709882e-21, -1.003089e-36, 2.569961e-21, -7.709882e-21, 
    1.027984e-20, 5.139921e-21, 1.28498e-20, -1.003089e-36, -1.003089e-36, 
    2.569961e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, -7.709882e-21, 
    -2.055969e-20, 0, 1.003089e-36, 5.139921e-21, -1.28498e-20, 
    -1.003089e-36, 2.569961e-21, 1.027984e-20, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 1.28498e-20, -7.709882e-21, -1.027984e-20, 5.139921e-21, 
    1.027984e-20, -2.569961e-21, 2.569961e-21, 5.139921e-21, 0, 
    -1.541976e-20, -1.541976e-20, -2.826957e-20, 1.798972e-20, -2.569961e-21, 
    -1.798972e-20, 5.139921e-21, 2.569961e-21, 1.027984e-20, 1.28498e-20, 
    1.541976e-20, -2.569961e-21, -1.541976e-20, 0, -2.055969e-20, 
    5.139921e-21, 1.027984e-20, -1.003089e-36, -2.569961e-21, -5.139921e-21, 
    1.003089e-36, 0, 2.569961e-21, 5.139921e-21, -2.569961e-21, 
    -5.139921e-21, 1.798972e-20, 2.055969e-20, 1.28498e-20, 2.569961e-21, 
    -1.541976e-20, 1.003089e-36, 2.569961e-21, -1.027984e-20, 5.139921e-21, 
    -1.027984e-20, -5.139921e-21, 7.709882e-21, 1.28498e-20, -1.28498e-20, 
    -1.28498e-20, -5.139921e-21, 1.541976e-20, -5.139921e-21, 7.709882e-21, 
    1.003089e-36, 1.541976e-20, 7.709882e-21, -2.569961e-21, -1.798972e-20, 
    2.569961e-21, 1.027984e-20, 2.569961e-21, -1.027984e-20, 1.003089e-36, 
    5.139921e-21, -1.798972e-20, -2.055969e-20, 1.28498e-20, 1.027984e-20, 
    2.569961e-21, 1.28498e-20, 1.003089e-36, -2.569961e-21, 2.569961e-21, 
    5.139921e-21, -1.027984e-20, -1.003089e-36, 5.139921e-21, -1.28498e-20, 
    1.28498e-20, -1.027984e-20, -1.798972e-20, -2.569961e-20, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, -2.055969e-20, 1.027984e-20, 
    2.569961e-21, 1.027984e-20, 7.709882e-21, 5.139921e-21, -1.28498e-20, 
    5.139921e-21, 1.027984e-20, -5.139921e-21, -5.015443e-37, -7.709882e-21,
  2.569961e-21, -7.709882e-21, -2.569961e-21, 0, -1.541976e-20, 
    -7.709882e-21, -2.569961e-21, 5.139921e-21, 7.709882e-21, 1.541976e-20, 
    5.139921e-21, 7.709882e-21, 2.569961e-21, 2.569961e-21, -5.139921e-21, 
    -7.709882e-21, 1.541976e-20, 1.003089e-36, -1.003089e-36, -7.709882e-21, 
    0, -7.709882e-21, -2.569961e-21, -1.28498e-20, -5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 2.569961e-21, 7.709882e-21, 7.709882e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, -7.709882e-21, -1.28498e-20, 
    -5.139921e-21, -7.709882e-21, 2.569961e-21, 1.027984e-20, 7.709882e-21, 
    -2.569961e-21, 2.569961e-21, 5.139921e-21, -5.139921e-21, 7.709882e-21, 
    1.027984e-20, 7.709882e-21, 1.28498e-20, 0, 1.027984e-20, 2.569961e-21, 
    1.027984e-20, 7.709882e-21, -1.28498e-20, -2.569961e-21, -5.139921e-21, 
    -7.709882e-21, -5.139921e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, 2.569961e-21, 1.003089e-36, -7.709882e-21, 0, 0, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, 0, 
    -7.709882e-21, -5.139921e-21, -5.139921e-21, 5.139921e-21, 1.027984e-20, 
    2.569961e-21, 5.139921e-21, -5.139921e-21, 2.569961e-21, 1.003089e-36, 0, 
    5.139921e-21, 2.569961e-21, -5.139921e-21, 2.569961e-21, -1.027984e-20, 
    -7.709882e-21, 5.139921e-21, 0, 1.28498e-20, 7.709882e-21, 1.027984e-20, 
    1.541976e-20, 2.569961e-21, 5.139921e-21, -1.003089e-36, -1.027984e-20, 
    -7.709882e-21, 0, -7.709882e-21, -2.569961e-21, -1.541976e-20, 
    -1.541976e-20, 2.569961e-21, 1.28498e-20, 2.569961e-21, 7.709882e-21, 
    -1.027984e-20, 1.003089e-36, -1.541976e-20, 5.139921e-21, 5.139921e-21, 
    -1.027984e-20, 1.027984e-20, -5.139921e-21, -1.798972e-20, -5.139921e-21, 
    5.139921e-21, -5.139921e-21, 2.569961e-21, -2.569961e-21, -1.027984e-20, 
    -2.569961e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, -5.139921e-21, 
    2.569961e-21, 7.709882e-21, 2.569961e-21, -1.798972e-20, -2.569961e-21, 
    -1.027984e-20, -5.139921e-21, 5.139921e-21, 1.003089e-36, 7.709882e-21, 
    5.139921e-21, 0, -1.027984e-20, 5.139921e-21, -1.541976e-20, 
    -1.541976e-20, 7.709882e-21, 5.139921e-21, -5.139921e-21, -1.541976e-20, 
    -5.139921e-21, 1.027984e-20, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -1.003089e-36, 5.139921e-21, -2.569961e-21, 5.139921e-21, 0, 
    -5.139921e-21, 1.027984e-20, 5.139921e-21, -1.027984e-20, -1.003089e-36, 
    -1.003089e-36, -2.055969e-20, 0, 5.139921e-21, -1.003089e-36, 
    -2.569961e-21, -5.139921e-21, -2.569961e-21, 0, -2.569961e-21, 
    2.569961e-21, -2.569961e-21, 0, -7.709882e-21, 0, -5.139921e-21, 
    -1.003089e-36, 5.139921e-21, -5.139921e-21, 1.003089e-36, -1.003089e-36, 
    7.709882e-21, 5.139921e-21, -5.139921e-21, -1.798972e-20, 1.003089e-36, 
    -2.569961e-21, 0, -7.709882e-21, -5.139921e-21, -7.709882e-21, 
    5.139921e-21, -1.28498e-20, -7.709882e-21, -7.709882e-21, -5.139921e-21, 
    5.139921e-21, -7.709882e-21, 2.569961e-21, 5.139921e-21, 2.569961e-21, 
    -7.709882e-21, 2.569961e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, 
    1.027984e-20, -2.569961e-21, 5.139921e-21, 2.569961e-21, 1.28498e-20, 
    2.569961e-21, 1.003089e-36, 7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -1.027984e-20, 7.709882e-21, 2.569961e-21, 0, 1.003089e-36, 5.139921e-21, 
    -7.709882e-21, -5.139921e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, 
    -5.139921e-21, -2.569961e-21, 1.28498e-20, 1.027984e-20, -1.003089e-36, 
    7.709882e-21, 1.027984e-20, 7.709882e-21, 2.569961e-21, -2.569961e-21, 
    -1.003089e-36, -5.139921e-21, -2.569961e-21, 7.709882e-21, 2.569961e-21, 
    7.709882e-21, -2.569961e-21, 7.709882e-21, -5.139921e-21, 5.139921e-21, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, 0, -1.027984e-20, 
    -1.28498e-20, 7.709882e-21, 1.027984e-20, -5.139921e-21, 2.312965e-20, 
    -5.139921e-21, 2.569961e-21, -1.003089e-36, 1.003089e-36, 2.569961e-21, 
    1.027984e-20, 7.709882e-21, -1.003089e-36, -2.569961e-21, 2.569961e-21, 
    1.027984e-20, -2.569961e-21, 5.139921e-21, -7.709882e-21, -7.709882e-21, 
    -2.569961e-21, 1.027984e-20, -7.709882e-21, 2.569961e-21, 7.709882e-21, 
    -1.003089e-36, 1.027984e-20, 0, -2.569961e-21, 1.541976e-20, 
    -2.569961e-21, 5.139921e-21, -1.541976e-20, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, 1.541976e-20, 7.709882e-21, -7.709882e-21, 5.139921e-21, 
    -7.709882e-21, 5.139921e-21, 0, 1.003089e-36, 1.003089e-36, 2.569961e-21, 
    2.569961e-21, -5.139921e-21, 7.709882e-21, 5.139921e-21, -2.569961e-21, 
    1.027984e-20, 5.139921e-21, 1.027984e-20, 0, 2.569961e-21, -7.709882e-21, 
    -2.569961e-21, -1.28498e-20, 7.709882e-21, 0, 2.569961e-21, 
    -2.569961e-21, 0, 1.541976e-20, 5.139921e-21, -1.541976e-20, 
    2.569961e-21, 1.027984e-20, -2.569961e-21, 7.709882e-21, 1.027984e-20, 
    2.569961e-21, -7.709882e-21, 0, 0, 5.139921e-21, -7.709882e-21, 
    5.139921e-21, -5.139921e-21, 2.055969e-20, -2.569961e-21,
  0, -7.709882e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, 0, 
    -2.569961e-21, -2.569961e-21, -2.569961e-21, -7.709882e-21, 
    -5.139921e-21, 7.709882e-21, -1.003089e-36, 2.569961e-21, 2.569961e-21, 
    -1.541976e-20, 5.139921e-21, 5.139921e-21, 7.709882e-21, -2.569961e-21, 
    0, -1.28498e-20, 1.28498e-20, -1.027984e-20, -1.003089e-36, 0, 
    -5.139921e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, -2.055969e-20, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, -5.139921e-21, -2.569961e-21, 
    7.709882e-21, -7.709882e-21, -2.569961e-21, -2.569961e-21, -5.139921e-21, 
    1.798972e-20, 2.569961e-21, 7.709882e-21, -2.569961e-21, 1.027984e-20, 
    -1.027984e-20, -5.139921e-21, 7.709882e-21, 7.709882e-21, 7.709882e-21, 
    -7.709882e-21, 7.709882e-21, 7.709882e-21, 7.709882e-21, -1.027984e-20, 
    5.139921e-21, 1.003089e-36, 2.569961e-21, -1.28498e-20, 2.569961e-21, 
    -7.709882e-21, -7.709882e-21, -2.569961e-21, 5.139921e-21, -7.709882e-21, 
    1.798972e-20, -2.826957e-20, 2.569961e-21, -2.569961e-21, 2.569961e-21, 
    5.139921e-21, -1.541976e-20, 2.569961e-21, 1.027984e-20, 7.709882e-21, 
    -1.027984e-20, -1.28498e-20, -1.027984e-20, -1.003089e-36, 5.139921e-21, 
    0, -1.027984e-20, -2.569961e-21, 2.569961e-21, 1.541976e-20, 
    -1.541976e-20, -2.569961e-21, 7.709882e-21, -2.569961e-21, -1.027984e-20, 
    2.569961e-21, -1.027984e-20, -2.569961e-21, -2.569961e-21, -1.28498e-20, 
    0, -7.709882e-21, -1.28498e-20, -1.003089e-36, 0, 1.027984e-20, 
    1.003089e-36, -5.139921e-21, -7.709882e-21, -7.709882e-21, 2.569961e-21, 
    7.709882e-21, 2.569961e-21, -7.709882e-21, -2.569961e-21, -5.139921e-21, 
    -5.139921e-21, -2.569961e-21, 1.003089e-36, 0, 7.709882e-21, 
    -1.28498e-20, -5.139921e-21, 1.027984e-20, 2.569961e-21, -7.709882e-21, 
    -5.139921e-21, 5.139921e-21, 0, -2.569961e-21, 7.709882e-21, 
    1.798972e-20, 1.28498e-20, -7.709882e-21, -2.569961e-21, 5.139921e-21, 
    -5.139921e-21, 0, 2.569961e-21, -7.709882e-21, 7.709882e-21, 
    -2.569961e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, -2.569961e-21, -7.709882e-21, -1.28498e-20, -1.28498e-20, 
    2.569961e-21, 5.139921e-21, -1.28498e-20, -7.709882e-21, -7.709882e-21, 
    -5.139921e-21, -2.569961e-21, 1.798972e-20, 1.28498e-20, -7.709882e-21, 
    -2.569961e-21, -5.139921e-21, -1.003089e-36, -2.055969e-20, 
    -2.569961e-21, 7.709882e-21, 1.027984e-20, 1.027984e-20, 7.709882e-21, 
    -1.28498e-20, -2.826957e-20, -2.569961e-21, -5.139921e-21, 1.541976e-20, 
    1.28498e-20, 7.709882e-21, -5.139921e-21, 1.027984e-20, 0, 7.709882e-21, 
    2.569961e-21, -2.569961e-21, 5.139921e-21, -5.139921e-21, 2.569961e-21, 
    1.027984e-20, -2.569961e-21, 7.709882e-21, 1.027984e-20, -1.003089e-36, 
    -5.139921e-21, -1.541976e-20, 0, 5.139921e-21, -1.28498e-20, 
    2.055969e-20, -2.569961e-21, -2.569961e-21, -1.798972e-20, -1.541976e-20, 
    0, 1.027984e-20, -2.569961e-21, 1.28498e-20, -1.027984e-20, 2.569961e-21, 
    5.139921e-21, -5.139921e-21, 1.027984e-20, 5.139921e-21, 5.139921e-21, 
    5.139921e-21, 2.055969e-20, 2.569961e-21, 1.28498e-20, -2.569961e-21, 
    -5.139921e-21, -1.28498e-20, 1.28498e-20, 2.569961e-21, -5.139921e-21, 
    2.569961e-21, -5.139921e-21, 0, -5.139921e-21, 2.569961e-21, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, -1.027984e-20, -5.139921e-21, 
    -2.569961e-21, 0, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, -7.709882e-21, -2.569961e-21, 5.139921e-21, 1.541976e-20, 
    -1.28498e-20, -1.798972e-20, -1.027984e-20, 7.709882e-21, -5.139921e-21, 
    1.027984e-20, 1.027984e-20, 0, -1.798972e-20, 7.709882e-21, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, 1.28498e-20, 5.139921e-21, 
    -1.003089e-36, 5.139921e-21, 2.569961e-21, 1.28498e-20, -1.003089e-36, 
    2.569961e-21, 5.139921e-21, -5.139921e-21, 7.709882e-21, -5.139921e-21, 
    2.569961e-21, 2.569961e-21, -7.709882e-21, -5.139921e-21, -7.709882e-21, 
    2.569961e-21, 7.709882e-21, 7.709882e-21, 2.569961e-21, -5.139921e-21, 
    2.569961e-21, 2.569961e-21, 2.569961e-21, -1.28498e-20, -1.027984e-20, 
    -1.28498e-20, -5.139921e-21, 0, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 7.709882e-21, -1.003089e-36, -1.003089e-36, 0, 
    -2.569961e-21, 1.28498e-20, 7.709882e-21, 7.709882e-21, -1.28498e-20, 
    2.569961e-21, 1.28498e-20, -2.569961e-21, -1.003089e-36, 7.709882e-21, 0, 
    7.709882e-21, 1.027984e-20, 1.003089e-36, -2.569961e-21, 1.28498e-20, 
    -1.541976e-20, -5.139921e-21, 1.003089e-36, 0, 5.139921e-21, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, 5.139921e-21, -2.569961e-21, 
    -2.569961e-21, -1.027984e-20, 5.139921e-21, 2.569961e-21, 1.003089e-36, 
    -1.28498e-20, 1.798972e-20, -2.055969e-20, -2.569961e-21, 0, 0, 
    1.027984e-20, 5.139921e-21, -7.709882e-21, 5.139921e-21, -2.569961e-21, 
    -1.798972e-20, 1.28498e-20, 5.139921e-21, 1.798972e-20, -1.798972e-20, 
    2.569961e-21, 2.569961e-21, 7.709882e-21,
  -1.027984e-20, -7.709882e-21, 1.28498e-20, -5.139921e-21, -5.139921e-21, 
    -1.003089e-36, -1.027984e-20, -1.28498e-20, -2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -1.798972e-20, 7.709882e-21, 7.709882e-21, 0, 
    2.569961e-21, -1.28498e-20, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -1.027984e-20, -5.139921e-21, 
    -2.569961e-20, -2.569961e-21, 7.709882e-21, 1.541976e-20, -2.569961e-21, 
    0, 0, 1.027984e-20, -5.139921e-21, -1.28498e-20, -1.541976e-20, 
    -1.541976e-20, 5.139921e-21, -2.569961e-21, 1.027984e-20, 2.055969e-20, 
    5.139921e-21, -7.709882e-21, -1.28498e-20, -7.709882e-21, 1.28498e-20, 
    2.569961e-21, 1.541976e-20, -2.569961e-21, -1.541976e-20, -5.139921e-21, 
    7.709882e-21, 2.569961e-21, 5.139921e-21, -2.569961e-21, -1.027984e-20, 
    1.28498e-20, -2.569961e-21, -1.798972e-20, 1.027984e-20, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, 7.709882e-21, -1.003089e-36, 5.139921e-21, 
    -5.139921e-21, -1.28498e-20, -5.139921e-21, -1.541976e-20, -1.027984e-20, 
    7.709882e-21, 3.340949e-20, 1.541976e-20, -1.027984e-20, 7.709882e-21, 
    1.541976e-20, 7.709882e-21, 5.139921e-21, -7.709882e-21, -5.139921e-21, 
    2.569961e-21, -1.541976e-20, -7.709882e-21, 1.003089e-36, -1.798972e-20, 
    1.28498e-20, -1.027984e-20, -7.709882e-21, 1.027984e-20, -1.541976e-20, 
    -1.027984e-20, -1.027984e-20, -2.569961e-21, -7.709882e-21, 1.027984e-20, 
    -1.28498e-20, 7.709882e-21, -1.28498e-20, 5.139921e-21, -1.28498e-20, 0, 
    2.569961e-21, 5.139921e-21, 1.027984e-20, 5.139921e-21, -5.139921e-21, 
    5.139921e-21, 2.569961e-21, -1.027984e-20, 1.027984e-20, 5.139921e-21, 
    -1.541976e-20, 1.28498e-20, -2.569961e-21, 5.139921e-21, -7.709882e-21, 
    -1.027984e-20, 2.569961e-21, 1.027984e-20, -2.569961e-21, 5.139921e-21, 
    1.003089e-36, -2.569961e-21, -5.139921e-21, 2.569961e-21, -5.139921e-21, 
    -1.003089e-36, 5.139921e-21, 2.569961e-21, -7.709882e-21, -7.709882e-21, 
    -5.139921e-21, 1.027984e-20, -5.139921e-21, 5.139921e-21, 1.003089e-36, 
    1.027984e-20, 7.709882e-21, 2.569961e-21, -5.139921e-21, 5.139921e-21, 
    -2.569961e-21, 1.003089e-36, 7.709882e-21, 2.569961e-21, -1.798972e-20, 
    -1.003089e-36, 7.709882e-21, 2.569961e-21, 7.709882e-21, 2.055969e-20, 
    -7.709882e-21, 7.709882e-21, 7.709882e-21, -1.798972e-20, -1.027984e-20, 
    5.139921e-21, -2.569961e-21, 1.798972e-20, 1.003089e-36, -2.569961e-21, 
    -7.709882e-21, 5.139921e-21, 7.709882e-21, -1.28498e-20, 2.569961e-21, 
    -2.569961e-21, 1.541976e-20, -1.003089e-36, 7.709882e-21, -5.139921e-21, 
    -2.569961e-21, 7.709882e-21, -5.139921e-21, 7.709882e-21, 7.709882e-21, 
    2.569961e-21, -5.139921e-21, -1.28498e-20, -2.569961e-21, -1.28498e-20, 
    -1.003089e-36, -5.139921e-21, -1.28498e-20, -7.709882e-21, 1.003089e-36, 
    7.709882e-21, 7.709882e-21, 1.28498e-20, 1.027984e-20, 1.027984e-20, 
    2.569961e-21, 1.003089e-36, -2.569961e-21, -1.798972e-20, 1.027984e-20, 
    -2.569961e-21, 2.569961e-20, 5.139921e-21, 0, -5.139921e-21, 
    1.027984e-20, 0, -1.027984e-20, -5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 1.28498e-20, 7.709882e-21, 2.569961e-21, 1.027984e-20, 
    2.055969e-20, -1.541976e-20, 7.709882e-21, 5.139921e-21, -5.139921e-21, 
    -1.003089e-36, 2.569961e-21, -5.139921e-21, 1.28498e-20, -1.28498e-20, 
    5.139921e-21, 0, 2.569961e-21, 1.798972e-20, 1.28498e-20, 5.139921e-21, 
    -7.709882e-21, 1.003089e-36, -1.027984e-20, -1.027984e-20, 7.709882e-21, 
    -1.027984e-20, -5.139921e-21, -2.569961e-20, -1.027984e-20, 2.312965e-20, 
    5.139921e-21, 1.798972e-20, 1.027984e-20, -7.709882e-21, 5.139921e-21, 
    1.027984e-20, 0, -1.28498e-20, 1.541976e-20, -7.709882e-21, 5.139921e-21, 
    5.139921e-21, -1.28498e-20, -1.541976e-20, 1.027984e-20, -1.28498e-20, 
    -7.709882e-21, -7.709882e-21, 1.027984e-20, 5.139921e-21, 5.139921e-21, 
    2.055969e-20, -1.027984e-20, -7.709882e-21, 2.569961e-21, -1.798972e-20, 
    2.569961e-21, -1.003089e-36, -2.569961e-21, -1.003089e-36, -1.798972e-20, 
    -1.027984e-20, -1.027984e-20, 2.569961e-21, 7.709882e-21, -1.027984e-20, 
    -7.709882e-21, 0, -2.312965e-20, -2.569961e-20, 0, 7.709882e-21, 0, 
    2.055969e-20, 2.569961e-21, -1.003089e-36, 1.28498e-20, 2.569961e-21, 
    -7.709882e-21, 1.027984e-20, 1.541976e-20, 2.569961e-21, -1.027984e-20, 
    -1.798972e-20, -2.055969e-20, 1.541976e-20, 1.541976e-20, -1.003089e-36, 
    -2.569961e-21, 0, 2.569961e-21, 7.709882e-21, -5.139921e-21, 
    -1.027984e-20, -7.709882e-21, -1.28498e-20, 5.139921e-21, -7.709882e-21, 
    7.709882e-21, 2.569961e-21, 1.541976e-20, 5.139921e-21, -5.139921e-21, 
    -1.28498e-20, 1.003089e-36, 1.28498e-20, 7.709882e-21, 2.569961e-21, 
    5.139921e-21, 1.003089e-36, 5.139921e-21, -7.709882e-21, 7.709882e-21, 
    -2.569961e-21, 7.709882e-21, -7.709882e-21, 5.139921e-21, 1.027984e-20, 
    -1.003089e-36, 1.003089e-36, -5.139921e-21, -1.027984e-20, -5.139921e-21, 
    -2.569961e-21, 1.541976e-20, 1.027984e-20, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, -1.027984e-20, 1.541976e-20,
  -5.139921e-21, -2.569961e-21, -2.569961e-21, -7.709882e-21, -1.541976e-20, 
    5.139921e-21, 2.569961e-21, 1.027984e-20, 2.312965e-20, 2.569961e-21, 
    1.28498e-20, -7.709882e-21, 1.28498e-20, -5.139921e-21, -1.027984e-20, 
    -1.28498e-20, 2.569961e-21, 1.28498e-20, -7.709882e-21, 1.027984e-20, 
    -2.569961e-21, 5.139921e-21, -2.312965e-20, 5.139921e-21, 1.003089e-36, 
    1.798972e-20, -2.569961e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, 
    1.027984e-20, 2.312965e-20, 2.569961e-21, -1.28498e-20, 1.28498e-20, 
    1.003089e-36, -1.798972e-20, 0, 2.569961e-20, -5.139921e-21, 
    1.027984e-20, -1.541976e-20, -2.569961e-21, -5.139921e-21, 2.569961e-21, 
    -2.569961e-21, -5.139921e-21, 5.139921e-21, -2.569961e-21, 1.28498e-20, 
    -2.569961e-21, -2.569961e-21, -7.709882e-21, 5.139921e-21, 5.139921e-21, 
    7.709882e-21, -2.569961e-21, -2.569961e-21, -2.569961e-20, -2.569961e-21, 
    -2.569961e-21, 1.027984e-20, -5.139921e-21, 2.826957e-20, 0, 
    -1.798972e-20, 5.139921e-21, -1.027984e-20, -2.569961e-20, -2.569961e-21, 
    -1.027984e-20, 2.312965e-20, -1.003089e-36, 1.003089e-36, 5.139921e-21, 
    -1.541976e-20, 7.709882e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, 
    5.139921e-21, 5.139921e-21, 2.569961e-21, 7.709882e-21, 1.027984e-20, 
    -2.569961e-21, -2.312965e-20, -1.027984e-20, 2.569961e-21, 2.569961e-20, 
    2.569961e-21, -7.709882e-21, 1.027984e-20, 2.312965e-20, -1.28498e-20, 
    -1.28498e-20, -1.027984e-20, 7.709882e-21, -1.798972e-20, 2.569961e-21, 
    -2.569961e-21, 1.541976e-20, 2.569961e-21, -1.798972e-20, -1.027984e-20, 
    5.139921e-21, 2.055969e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    5.139921e-21, 2.569961e-21, 1.003089e-36, 0, -2.569961e-21, 1.28498e-20, 
    2.826957e-20, 1.003089e-36, 0, -1.541976e-20, 1.28498e-20, -7.709882e-21, 
    -1.798972e-20, 2.569961e-21, 2.055969e-20, -2.569961e-21, -2.569961e-21, 
    1.027984e-20, -2.569961e-20, -2.569961e-21, 1.798972e-20, -1.027984e-20, 
    1.027984e-20, 1.28498e-20, 2.569961e-21, 1.541976e-20, -1.28498e-20, 
    5.139921e-21, 1.28498e-20, -2.569961e-21, 1.027984e-20, 7.709882e-21, 
    1.541976e-20, -5.139921e-21, -2.312965e-20, 1.027984e-20, 2.569961e-21, 
    -1.027984e-20, 1.798972e-20, 1.027984e-20, -7.709882e-21, -1.027984e-20, 
    1.003089e-36, -7.709882e-21, -1.027984e-20, 2.569961e-20, 5.139921e-21, 
    2.569961e-21, 2.055969e-20, -2.569961e-21, 2.569961e-21, 2.055969e-20, 
    2.569961e-21, 1.027984e-20, -1.798972e-20, -1.28498e-20, 1.28498e-20, 
    -1.798972e-20, 0, -2.055969e-20, -1.027984e-20, 7.709882e-21, 
    -1.027984e-20, 1.28498e-20, -1.027984e-20, 1.28498e-20, -5.139921e-21, 
    7.709882e-21, 2.569961e-21, 1.28498e-20, 2.569961e-21, -2.569961e-21, 
    1.003089e-36, -2.569961e-21, 2.569961e-21, 7.709882e-21, 7.709882e-21, 
    -1.027984e-20, -5.139921e-21, -7.709882e-21, 7.709882e-21, -1.28498e-20, 
    1.027984e-20, 1.28498e-20, -2.569961e-21, -2.569961e-21, -1.027984e-20, 
    -1.027984e-20, -2.055969e-20, -1.541976e-20, 1.28498e-20, 1.28498e-20, 
    7.709882e-21, 7.709882e-21, -1.541976e-20, -1.541976e-20, -5.139921e-21, 
    -7.709882e-21, -1.798972e-20, -5.139921e-21, 5.139921e-21, -7.709882e-21, 
    -2.569961e-21, -7.709882e-21, -3.009266e-36, -1.027984e-20, 
    -2.312965e-20, 1.027984e-20, 1.003089e-36, 2.569961e-21, 1.798972e-20, 
    -1.28498e-20, -1.027984e-20, 7.709882e-21, 2.826957e-20, -1.28498e-20, 
    -5.139921e-21, -2.055969e-20, -7.709882e-21, -5.139921e-21, 
    -1.798972e-20, -5.139921e-21, -2.569961e-21, 1.28498e-20, -1.28498e-20, 
    -1.027984e-20, -1.027984e-20, 1.541976e-20, 2.569961e-21, -2.055969e-20, 
    1.28498e-20, -1.003089e-36, 2.569961e-21, -1.027984e-20, -2.569961e-21, 
    7.709882e-21, -2.569961e-21, 1.28498e-20, 5.139921e-21, -1.003089e-36, 
    2.569961e-21, 5.139921e-21, 2.569961e-21, -5.015443e-37, -1.798972e-20, 
    1.798972e-20, 7.709882e-21, -1.541976e-20, -1.003089e-36, -2.569961e-20, 
    -1.28498e-20, 5.139921e-21, -5.139921e-21, 1.28498e-20, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, -2.569961e-21, -5.139921e-21, 
    0, 1.541976e-20, -5.139921e-21, 1.003089e-36, 1.28498e-20, 5.139921e-21, 
    -2.312965e-20, 1.003089e-36, -1.541976e-20, -7.709882e-21, -1.027984e-20, 
    -1.027984e-20, 5.139921e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, 
    1.798972e-20, -7.709882e-21, 2.569961e-21, -2.569961e-20, -1.027984e-20, 
    -1.003089e-36, -1.027984e-20, 2.569961e-21, -2.312965e-20, 1.027984e-20, 
    2.569961e-21, -5.139921e-21, -5.139921e-21, 2.569961e-21, 5.139921e-21, 
    1.027984e-20, -7.709882e-21, 1.541976e-20, -1.027984e-20, 2.569961e-21, 
    7.709882e-21, 1.027984e-20, -7.709882e-21, 5.139921e-21, 1.003089e-36, 
    -1.541976e-20, -7.709882e-21, -2.569961e-21, -1.003089e-36, 2.569961e-21, 
    -1.003089e-36, -7.709882e-21, 1.28498e-20, -1.003089e-36, -1.798972e-20, 
    -2.055969e-20, -7.709882e-21, -1.541976e-20, -1.027984e-20, 
    -2.569961e-21, -7.709882e-21, -1.027984e-20, -7.709882e-21, 2.569961e-21, 
    1.28498e-20, 2.569961e-21, 1.541976e-20, -1.28498e-20, -2.569961e-21, 
    1.541976e-20, -5.139921e-21, -5.139921e-21,
  6.259414e-29, 6.25942e-29, 6.259419e-29, 6.259424e-29, 6.259422e-29, 
    6.259425e-29, 6.259416e-29, 6.25942e-29, 6.259417e-29, 6.259414e-29, 
    6.259434e-29, 6.259425e-29, 6.259444e-29, 6.259438e-29, 6.259453e-29, 
    6.259443e-29, 6.259456e-29, 6.259453e-29, 6.259461e-29, 6.259459e-29, 
    6.259468e-29, 6.259462e-29, 6.259473e-29, 6.259466e-29, 6.259467e-29, 
    6.259461e-29, 6.259426e-29, 6.259433e-29, 6.259426e-29, 6.259427e-29, 
    6.259426e-29, 6.259422e-29, 6.259419e-29, 6.259414e-29, 6.259414e-29, 
    6.259419e-29, 6.259428e-29, 6.259425e-29, 6.259432e-29, 6.259432e-29, 
    6.25944e-29, 6.259437e-29, 6.259451e-29, 6.259447e-29, 6.259459e-29, 
    6.259456e-29, 6.259458e-29, 6.259458e-29, 6.259458e-29, 6.259454e-29, 
    6.259456e-29, 6.259452e-29, 6.259437e-29, 6.259441e-29, 6.259429e-29, 
    6.259421e-29, 6.259416e-29, 6.259412e-29, 6.259413e-29, 6.259413e-29, 
    6.259419e-29, 6.259423e-29, 6.259427e-29, 6.259429e-29, 6.259432e-29, 
    6.259439e-29, 6.259443e-29, 6.259452e-29, 6.25945e-29, 6.259453e-29, 
    6.259455e-29, 6.259459e-29, 6.259459e-29, 6.259461e-29, 6.259453e-29, 
    6.259458e-29, 6.259449e-29, 6.259452e-29, 6.259432e-29, 6.259425e-29, 
    6.259422e-29, 6.259419e-29, 6.259413e-29, 6.259417e-29, 6.259416e-29, 
    6.25942e-29, 6.259423e-29, 6.259421e-29, 6.259429e-29, 6.259426e-29, 
    6.259443e-29, 6.259436e-29, 6.259455e-29, 6.25945e-29, 6.259456e-29, 
    6.259453e-29, 6.259458e-29, 6.259454e-29, 6.259461e-29, 6.259463e-29, 
    6.259462e-29, 6.259467e-29, 6.259453e-29, 6.259458e-29, 6.259421e-29, 
    6.259422e-29, 6.259422e-29, 6.259418e-29, 6.259417e-29, 6.259414e-29, 
    6.259417e-29, 6.259419e-29, 6.259423e-29, 6.259425e-29, 6.259427e-29, 
    6.259432e-29, 6.259438e-29, 6.259445e-29, 6.259451e-29, 6.259455e-29, 
    6.259452e-29, 6.259454e-29, 6.259452e-29, 6.259451e-29, 6.259463e-29, 
    6.259456e-29, 6.259466e-29, 6.259466e-29, 6.259461e-29, 6.259466e-29, 
    6.259422e-29, 6.25942e-29, 6.259416e-29, 6.259419e-29, 6.259413e-29, 
    6.259417e-29, 6.259419e-29, 6.259426e-29, 6.259428e-29, 6.259429e-29, 
    6.259433e-29, 6.259437e-29, 6.259444e-29, 6.25945e-29, 6.259455e-29, 
    6.259455e-29, 6.259455e-29, 6.259456e-29, 6.259453e-29, 6.259457e-29, 
    6.259458e-29, 6.259456e-29, 6.259466e-29, 6.259463e-29, 6.259466e-29, 
    6.259464e-29, 6.259421e-29, 6.259423e-29, 6.259422e-29, 6.259424e-29, 
    6.259422e-29, 6.259429e-29, 6.259431e-29, 6.259441e-29, 6.259437e-29, 
    6.259443e-29, 6.259437e-29, 6.259438e-29, 6.259443e-29, 6.259438e-29, 
    6.25945e-29, 6.259441e-29, 6.259456e-29, 6.259449e-29, 6.259457e-29, 
    6.259455e-29, 6.259458e-29, 6.259461e-29, 6.259463e-29, 6.259469e-29, 
    6.259467e-29, 6.259472e-29, 6.259426e-29, 6.259429e-29, 6.259428e-29, 
    6.259431e-29, 6.259434e-29, 6.259438e-29, 6.259446e-29, 6.259443e-29, 
    6.259448e-29, 6.259449e-29, 6.259441e-29, 6.259446e-29, 6.259431e-29, 
    6.259433e-29, 6.259432e-29, 6.259426e-29, 6.259443e-29, 6.259435e-29, 
    6.259451e-29, 6.259446e-29, 6.25946e-29, 6.259453e-29, 6.259467e-29, 
    6.259473e-29, 6.259478e-29, 6.259485e-29, 6.25943e-29, 6.259428e-29, 
    6.259432e-29, 6.259437e-29, 6.259441e-29, 6.259446e-29, 6.259447e-29, 
    6.259448e-29, 6.259451e-29, 6.259453e-29, 6.259449e-29, 6.259454e-29, 
    6.259434e-29, 6.259444e-29, 6.259428e-29, 6.259432e-29, 6.259436e-29, 
    6.259435e-29, 6.259443e-29, 6.259444e-29, 6.259452e-29, 6.259448e-29, 
    6.259472e-29, 6.259461e-29, 6.25949e-29, 6.259482e-29, 6.259428e-29, 
    6.25943e-29, 6.259439e-29, 6.259435e-29, 6.259447e-29, 6.25945e-29, 
    6.259452e-29, 6.259455e-29, 6.259455e-29, 6.259457e-29, 6.259455e-29, 
    6.259457e-29, 6.259446e-29, 6.259451e-29, 6.259438e-29, 6.259441e-29, 
    6.25944e-29, 6.259438e-29, 6.259443e-29, 6.259449e-29, 6.259449e-29, 
    6.25945e-29, 6.259455e-29, 6.259447e-29, 6.259473e-29, 6.259456e-29, 
    6.259433e-29, 6.259438e-29, 6.259438e-29, 6.259437e-29, 6.259449e-29, 
    6.259445e-29, 6.259457e-29, 6.259454e-29, 6.259459e-29, 6.259456e-29, 
    6.259456e-29, 6.259453e-29, 6.25945e-29, 6.259445e-29, 6.25944e-29, 
    6.259437e-29, 6.259438e-29, 6.259441e-29, 6.259449e-29, 6.259455e-29, 
    6.259454e-29, 6.259459e-29, 6.259446e-29, 6.259452e-29, 6.259449e-29, 
    6.259455e-29, 6.259443e-29, 6.259453e-29, 6.25944e-29, 6.259441e-29, 
    6.259444e-29, 6.259452e-29, 6.259453e-29, 6.259455e-29, 6.259454e-29, 
    6.259449e-29, 6.259448e-29, 6.259444e-29, 6.259444e-29, 6.259441e-29, 
    6.259438e-29, 6.259441e-29, 6.259443e-29, 6.259449e-29, 6.259455e-29, 
    6.259461e-29, 6.259462e-29, 6.259469e-29, 6.259463e-29, 6.259473e-29, 
    6.259465e-29, 6.259479e-29, 6.259453e-29, 6.259464e-29, 6.259445e-29, 
    6.259447e-29, 6.259451e-29, 6.259459e-29, 6.259455e-29, 6.25946e-29, 
    6.259448e-29, 6.259442e-29, 6.25944e-29, 6.259437e-29, 6.25944e-29, 
    6.25944e-29, 6.259443e-29, 6.259442e-29, 6.259449e-29, 6.259446e-29, 
    6.259456e-29, 6.25946e-29, 6.259472e-29, 6.259479e-29, 6.259485e-29, 
    6.259489e-29, 6.25949e-29, 6.25949e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N_TO_SOIL1N =
  2.19423e-10, 2.203886e-10, 2.202009e-10, 2.209797e-10, 2.205476e-10, 
    2.210576e-10, 2.196188e-10, 2.204269e-10, 2.19911e-10, 2.195099e-10, 
    2.22491e-10, 2.210144e-10, 2.240248e-10, 2.23083e-10, 2.254486e-10, 
    2.238782e-10, 2.257653e-10, 2.254033e-10, 2.264927e-10, 2.261806e-10, 
    2.275741e-10, 2.266368e-10, 2.282964e-10, 2.273502e-10, 2.274983e-10, 
    2.266058e-10, 2.213115e-10, 2.223072e-10, 2.212525e-10, 2.213945e-10, 
    2.213308e-10, 2.205566e-10, 2.201664e-10, 2.193492e-10, 2.194976e-10, 
    2.200978e-10, 2.214584e-10, 2.209965e-10, 2.221605e-10, 2.221342e-10, 
    2.234301e-10, 2.228458e-10, 2.250238e-10, 2.244048e-10, 2.261936e-10, 
    2.257438e-10, 2.261725e-10, 2.260425e-10, 2.261742e-10, 2.255144e-10, 
    2.257971e-10, 2.252165e-10, 2.229552e-10, 2.236198e-10, 2.216377e-10, 
    2.204459e-10, 2.196542e-10, 2.190924e-10, 2.191719e-10, 2.193233e-10, 
    2.201013e-10, 2.208327e-10, 2.213902e-10, 2.21763e-10, 2.221304e-10, 
    2.232426e-10, 2.238311e-10, 2.25149e-10, 2.249112e-10, 2.253141e-10, 
    2.25699e-10, 2.263453e-10, 2.262389e-10, 2.265236e-10, 2.253035e-10, 
    2.261144e-10, 2.247757e-10, 2.251418e-10, 2.222304e-10, 2.211211e-10, 
    2.206497e-10, 2.202369e-10, 2.192329e-10, 2.199263e-10, 2.19653e-10, 
    2.203032e-10, 2.207164e-10, 2.20512e-10, 2.217732e-10, 2.212829e-10, 
    2.23866e-10, 2.227534e-10, 2.256541e-10, 2.2496e-10, 2.258205e-10, 
    2.253814e-10, 2.261338e-10, 2.254566e-10, 2.266296e-10, 2.26885e-10, 
    2.267105e-10, 2.273809e-10, 2.254191e-10, 2.261725e-10, 2.205063e-10, 
    2.205396e-10, 2.206949e-10, 2.200124e-10, 2.199706e-10, 2.193451e-10, 
    2.199017e-10, 2.201387e-10, 2.207403e-10, 2.210962e-10, 2.214345e-10, 
    2.221783e-10, 2.23009e-10, 2.241705e-10, 2.25005e-10, 2.255644e-10, 
    2.252214e-10, 2.255242e-10, 2.251857e-10, 2.25027e-10, 2.267893e-10, 
    2.257998e-10, 2.272845e-10, 2.272023e-10, 2.265304e-10, 2.272116e-10, 
    2.20563e-10, 2.203712e-10, 2.197054e-10, 2.202265e-10, 2.19277e-10, 
    2.198085e-10, 2.201141e-10, 2.212932e-10, 2.215522e-10, 2.217924e-10, 
    2.222669e-10, 2.228757e-10, 2.239438e-10, 2.248731e-10, 2.257214e-10, 
    2.256593e-10, 2.256811e-10, 2.258707e-10, 2.254012e-10, 2.259477e-10, 
    2.260395e-10, 2.257996e-10, 2.271913e-10, 2.267937e-10, 2.272006e-10, 
    2.269417e-10, 2.204336e-10, 2.207563e-10, 2.205819e-10, 2.209098e-10, 
    2.206788e-10, 2.217061e-10, 2.220141e-10, 2.234552e-10, 2.228637e-10, 
    2.23805e-10, 2.229593e-10, 2.231092e-10, 2.238358e-10, 2.23005e-10, 
    2.248219e-10, 2.235902e-10, 2.25878e-10, 2.246481e-10, 2.259551e-10, 
    2.257177e-10, 2.261107e-10, 2.264627e-10, 2.269055e-10, 2.277225e-10, 
    2.275333e-10, 2.282165e-10, 2.212374e-10, 2.21656e-10, 2.216191e-10, 
    2.220572e-10, 2.223811e-10, 2.230833e-10, 2.242094e-10, 2.237859e-10, 
    2.245634e-10, 2.247195e-10, 2.235383e-10, 2.242635e-10, 2.219361e-10, 
    2.223122e-10, 2.220883e-10, 2.212704e-10, 2.238836e-10, 2.225425e-10, 
    2.250188e-10, 2.242923e-10, 2.264125e-10, 2.253581e-10, 2.274291e-10, 
    2.283145e-10, 2.291477e-10, 2.301215e-10, 2.218844e-10, 2.216e-10, 
    2.221092e-10, 2.228139e-10, 2.234676e-10, 2.243366e-10, 2.244255e-10, 
    2.245884e-10, 2.250101e-10, 2.253647e-10, 2.246399e-10, 2.254536e-10, 
    2.223994e-10, 2.239999e-10, 2.214925e-10, 2.222476e-10, 2.227723e-10, 
    2.225421e-10, 2.237375e-10, 2.240193e-10, 2.251642e-10, 2.245723e-10, 
    2.28096e-10, 2.265371e-10, 2.308629e-10, 2.296541e-10, 2.215006e-10, 
    2.218834e-10, 2.232157e-10, 2.225818e-10, 2.243946e-10, 2.248409e-10, 
    2.252036e-10, 2.256673e-10, 2.257174e-10, 2.259921e-10, 2.255419e-10, 
    2.259743e-10, 2.243385e-10, 2.250695e-10, 2.230634e-10, 2.235517e-10, 
    2.233271e-10, 2.230807e-10, 2.238411e-10, 2.246513e-10, 2.246686e-10, 
    2.249283e-10, 2.256604e-10, 2.24402e-10, 2.282973e-10, 2.258917e-10, 
    2.223009e-10, 2.230382e-10, 2.231435e-10, 2.228579e-10, 2.247961e-10, 
    2.240938e-10, 2.259854e-10, 2.254742e-10, 2.263118e-10, 2.258956e-10, 
    2.258343e-10, 2.252997e-10, 2.249669e-10, 2.241261e-10, 2.234419e-10, 
    2.228993e-10, 2.230255e-10, 2.236215e-10, 2.247008e-10, 2.257219e-10, 
    2.254982e-10, 2.262481e-10, 2.242632e-10, 2.250955e-10, 2.247739e-10, 
    2.256126e-10, 2.237747e-10, 2.253399e-10, 2.233746e-10, 2.235469e-10, 
    2.240799e-10, 2.25152e-10, 2.253892e-10, 2.256424e-10, 2.254861e-10, 
    2.247282e-10, 2.24604e-10, 2.240669e-10, 2.239187e-10, 2.235094e-10, 
    2.231706e-10, 2.234802e-10, 2.238053e-10, 2.247285e-10, 2.255606e-10, 
    2.264677e-10, 2.266897e-10, 2.277497e-10, 2.268868e-10, 2.283107e-10, 
    2.271002e-10, 2.291956e-10, 2.254305e-10, 2.270646e-10, 2.241041e-10, 
    2.244231e-10, 2.249999e-10, 2.26323e-10, 2.256087e-10, 2.264441e-10, 
    2.245992e-10, 2.23642e-10, 2.233943e-10, 2.229323e-10, 2.234049e-10, 
    2.233665e-10, 2.238187e-10, 2.236734e-10, 2.247592e-10, 2.241759e-10, 
    2.258328e-10, 2.264375e-10, 2.281449e-10, 2.291917e-10, 2.302572e-10, 
    2.307276e-10, 2.308707e-10, 2.309306e-10 ;

 SOIL2N_TO_SOIL3N =
  1.567307e-11, 1.574204e-11, 1.572863e-11, 1.578426e-11, 1.57534e-11, 
    1.578983e-11, 1.568705e-11, 1.574478e-11, 1.570793e-11, 1.567928e-11, 
    1.589222e-11, 1.578674e-11, 1.600177e-11, 1.59345e-11, 1.610347e-11, 
    1.59913e-11, 1.612609e-11, 1.610024e-11, 1.617805e-11, 1.615576e-11, 
    1.625529e-11, 1.618834e-11, 1.630688e-11, 1.62393e-11, 1.624987e-11, 
    1.618613e-11, 1.580797e-11, 1.587909e-11, 1.580375e-11, 1.58139e-11, 
    1.580934e-11, 1.575404e-11, 1.572617e-11, 1.56678e-11, 1.56784e-11, 
    1.572127e-11, 1.581846e-11, 1.578546e-11, 1.586861e-11, 1.586673e-11, 
    1.595929e-11, 1.591756e-11, 1.607313e-11, 1.602892e-11, 1.615669e-11, 
    1.612455e-11, 1.615518e-11, 1.614589e-11, 1.61553e-11, 1.610817e-11, 
    1.612837e-11, 1.60869e-11, 1.592537e-11, 1.597284e-11, 1.583127e-11, 
    1.574614e-11, 1.568959e-11, 1.564946e-11, 1.565513e-11, 1.566595e-11, 
    1.572152e-11, 1.577377e-11, 1.581358e-11, 1.584022e-11, 1.586646e-11, 
    1.59459e-11, 1.598794e-11, 1.608207e-11, 1.606509e-11, 1.609387e-11, 
    1.612136e-11, 1.616752e-11, 1.615992e-11, 1.618026e-11, 1.60931e-11, 
    1.615103e-11, 1.605541e-11, 1.608156e-11, 1.58736e-11, 1.579436e-11, 
    1.576069e-11, 1.573121e-11, 1.565949e-11, 1.570902e-11, 1.56895e-11, 
    1.573594e-11, 1.576546e-11, 1.575086e-11, 1.584094e-11, 1.580592e-11, 
    1.599043e-11, 1.591096e-11, 1.611815e-11, 1.606857e-11, 1.613004e-11, 
    1.609867e-11, 1.615241e-11, 1.610405e-11, 1.618783e-11, 1.620607e-11, 
    1.619361e-11, 1.624149e-11, 1.610137e-11, 1.615518e-11, 1.575045e-11, 
    1.575283e-11, 1.576392e-11, 1.571517e-11, 1.571219e-11, 1.566751e-11, 
    1.570726e-11, 1.572419e-11, 1.576717e-11, 1.579259e-11, 1.581675e-11, 
    1.586988e-11, 1.592921e-11, 1.601218e-11, 1.607178e-11, 1.611174e-11, 
    1.608724e-11, 1.610887e-11, 1.608469e-11, 1.607336e-11, 1.619924e-11, 
    1.612855e-11, 1.623461e-11, 1.622874e-11, 1.618074e-11, 1.62294e-11, 
    1.57545e-11, 1.57408e-11, 1.569324e-11, 1.573046e-11, 1.566264e-11, 
    1.570061e-11, 1.572243e-11, 1.580666e-11, 1.582516e-11, 1.584232e-11, 
    1.58762e-11, 1.591969e-11, 1.599599e-11, 1.606236e-11, 1.612296e-11, 
    1.611852e-11, 1.612008e-11, 1.613362e-11, 1.610009e-11, 1.613912e-11, 
    1.614568e-11, 1.612854e-11, 1.622795e-11, 1.619955e-11, 1.622861e-11, 
    1.621012e-11, 1.574526e-11, 1.576831e-11, 1.575585e-11, 1.577927e-11, 
    1.576277e-11, 1.583615e-11, 1.585815e-11, 1.596108e-11, 1.591884e-11, 
    1.598607e-11, 1.592567e-11, 1.593637e-11, 1.598827e-11, 1.592893e-11, 
    1.60587e-11, 1.597072e-11, 1.613414e-11, 1.604629e-11, 1.613965e-11, 
    1.61227e-11, 1.615077e-11, 1.617591e-11, 1.620753e-11, 1.626589e-11, 
    1.625238e-11, 1.630118e-11, 1.580267e-11, 1.583257e-11, 1.582994e-11, 
    1.586123e-11, 1.588437e-11, 1.593452e-11, 1.601496e-11, 1.598471e-11, 
    1.604024e-11, 1.605139e-11, 1.596702e-11, 1.601882e-11, 1.585258e-11, 
    1.587944e-11, 1.586345e-11, 1.580503e-11, 1.599168e-11, 1.589589e-11, 
    1.607277e-11, 1.602088e-11, 1.617232e-11, 1.609701e-11, 1.624494e-11, 
    1.630818e-11, 1.63677e-11, 1.643725e-11, 1.584889e-11, 1.582857e-11, 
    1.586495e-11, 1.591527e-11, 1.596197e-11, 1.602404e-11, 1.60304e-11, 
    1.604203e-11, 1.607215e-11, 1.609748e-11, 1.60457e-11, 1.610382e-11, 
    1.588567e-11, 1.6e-11, 1.582089e-11, 1.587483e-11, 1.591231e-11, 
    1.589586e-11, 1.598125e-11, 1.600138e-11, 1.608316e-11, 1.604088e-11, 
    1.629257e-11, 1.618122e-11, 1.649021e-11, 1.640386e-11, 1.582147e-11, 
    1.584882e-11, 1.594398e-11, 1.58987e-11, 1.602819e-11, 1.606006e-11, 
    1.608597e-11, 1.611909e-11, 1.612267e-11, 1.614229e-11, 1.611013e-11, 
    1.614102e-11, 1.602418e-11, 1.607639e-11, 1.59331e-11, 1.596798e-11, 
    1.595193e-11, 1.593434e-11, 1.598865e-11, 1.604652e-11, 1.604776e-11, 
    1.606631e-11, 1.61186e-11, 1.602871e-11, 1.630695e-11, 1.613512e-11, 
    1.587863e-11, 1.59313e-11, 1.593882e-11, 1.591842e-11, 1.605687e-11, 
    1.60067e-11, 1.614182e-11, 1.61053e-11, 1.616513e-11, 1.61354e-11, 
    1.613102e-11, 1.609284e-11, 1.606907e-11, 1.6009e-11, 1.596013e-11, 
    1.592138e-11, 1.593039e-11, 1.597296e-11, 1.605006e-11, 1.612299e-11, 
    1.610702e-11, 1.616058e-11, 1.60188e-11, 1.607825e-11, 1.605528e-11, 
    1.611519e-11, 1.598391e-11, 1.609571e-11, 1.595533e-11, 1.596764e-11, 
    1.600571e-11, 1.608229e-11, 1.609923e-11, 1.611732e-11, 1.610615e-11, 
    1.605202e-11, 1.604315e-11, 1.600478e-11, 1.599419e-11, 1.596496e-11, 
    1.594076e-11, 1.596287e-11, 1.598609e-11, 1.605204e-11, 1.611147e-11, 
    1.617627e-11, 1.619212e-11, 1.626783e-11, 1.62062e-11, 1.630791e-11, 
    1.622144e-11, 1.637111e-11, 1.610218e-11, 1.62189e-11, 1.600744e-11, 
    1.603022e-11, 1.607143e-11, 1.616593e-11, 1.611491e-11, 1.617458e-11, 
    1.60428e-11, 1.597443e-11, 1.595674e-11, 1.592374e-11, 1.595749e-11, 
    1.595475e-11, 1.598705e-11, 1.597667e-11, 1.605423e-11, 1.601257e-11, 
    1.613091e-11, 1.61741e-11, 1.629607e-11, 1.637084e-11, 1.644694e-11, 
    1.648054e-11, 1.649077e-11, 1.649504e-11 ;

 SOIL2N_vr =
  1.818769, 1.818771, 1.81877, 1.818772, 1.818771, 1.818772, 1.81877, 
    1.818771, 1.81877, 1.818769, 1.818774, 1.818772, 1.818776, 1.818775, 
    1.818779, 1.818776, 1.818779, 1.818779, 1.81878, 1.81878, 1.818782, 
    1.818781, 1.818783, 1.818782, 1.818782, 1.818781, 1.818772, 1.818774, 
    1.818772, 1.818772, 1.818772, 1.818771, 1.81877, 1.818769, 1.818769, 
    1.81877, 1.818772, 1.818772, 1.818774, 1.818774, 1.818776, 1.818775, 
    1.818778, 1.818777, 1.81878, 1.818779, 1.81878, 1.81878, 1.81878, 
    1.818779, 1.818779, 1.818778, 1.818775, 1.818776, 1.818773, 1.818771, 
    1.81877, 1.818769, 1.818769, 1.818769, 1.81877, 1.818771, 1.818772, 
    1.818773, 1.818774, 1.818775, 1.818776, 1.818778, 1.818778, 1.818779, 
    1.818779, 1.81878, 1.81878, 1.81878, 1.818779, 1.81878, 1.818778, 
    1.818778, 1.818774, 1.818772, 1.818771, 1.818771, 1.818769, 1.81877, 
    1.81877, 1.818771, 1.818771, 1.818771, 1.818773, 1.818772, 1.818776, 
    1.818774, 1.818779, 1.818778, 1.818779, 1.818779, 1.81878, 1.818779, 
    1.818781, 1.818781, 1.818781, 1.818782, 1.818779, 1.81878, 1.818771, 
    1.818771, 1.818771, 1.81877, 1.81877, 1.818769, 1.81877, 1.81877, 
    1.818771, 1.818772, 1.818772, 1.818774, 1.818775, 1.818777, 1.818778, 
    1.818779, 1.818778, 1.818779, 1.818778, 1.818778, 1.818781, 1.818779, 
    1.818782, 1.818781, 1.81878, 1.818781, 1.818771, 1.818771, 1.81877, 
    1.818771, 1.818769, 1.81877, 1.81877, 1.818772, 1.818773, 1.818773, 
    1.818774, 1.818775, 1.818776, 1.818778, 1.818779, 1.818779, 1.818779, 
    1.818779, 1.818779, 1.81878, 1.81878, 1.818779, 1.818781, 1.818781, 
    1.818781, 1.818781, 1.818771, 1.818771, 1.818771, 1.818772, 1.818771, 
    1.818773, 1.818773, 1.818776, 1.818775, 1.818776, 1.818775, 1.818775, 
    1.818776, 1.818775, 1.818778, 1.818776, 1.818779, 1.818777, 1.81878, 
    1.818779, 1.81878, 1.81878, 1.818781, 1.818782, 1.818782, 1.818783, 
    1.818772, 1.818773, 1.818773, 1.818773, 1.818774, 1.818775, 1.818777, 
    1.818776, 1.818777, 1.818778, 1.818776, 1.818777, 1.818773, 1.818774, 
    1.818773, 1.818772, 1.818776, 1.818774, 1.818778, 1.818777, 1.81878, 
    1.818779, 1.818782, 1.818783, 1.818785, 1.818786, 1.818773, 1.818773, 
    1.818774, 1.818775, 1.818776, 1.818777, 1.818777, 1.818777, 1.818778, 
    1.818779, 1.818777, 1.818779, 1.818774, 1.818776, 1.818773, 1.818774, 
    1.818775, 1.818774, 1.818776, 1.818776, 1.818778, 1.818777, 1.818783, 
    1.81878, 1.818787, 1.818785, 1.818773, 1.818773, 1.818775, 1.818774, 
    1.818777, 1.818778, 1.818778, 1.818779, 1.818779, 1.81878, 1.818779, 
    1.81878, 1.818777, 1.818778, 1.818775, 1.818776, 1.818775, 1.818775, 
    1.818776, 1.818777, 1.818778, 1.818778, 1.818779, 1.818777, 1.818783, 
    1.818779, 1.818774, 1.818775, 1.818775, 1.818775, 1.818778, 1.818777, 
    1.81878, 1.818779, 1.81878, 1.818779, 1.818779, 1.818779, 1.818778, 
    1.818777, 1.818776, 1.818775, 1.818775, 1.818776, 1.818778, 1.818779, 
    1.818779, 1.81878, 1.818777, 1.818778, 1.818778, 1.818779, 1.818776, 
    1.818779, 1.818776, 1.818776, 1.818777, 1.818778, 1.818779, 1.818779, 
    1.818779, 1.818778, 1.818777, 1.818777, 1.818776, 1.818776, 1.818775, 
    1.818776, 1.818776, 1.818778, 1.818779, 1.81878, 1.818781, 1.818782, 
    1.818781, 1.818783, 1.818781, 1.818785, 1.818779, 1.818781, 1.818777, 
    1.818777, 1.818778, 1.81878, 1.818779, 1.81878, 1.818777, 1.818776, 
    1.818776, 1.818775, 1.818776, 1.818775, 1.818776, 1.818776, 1.818778, 
    1.818777, 1.818779, 1.81878, 1.818783, 1.818785, 1.818786, 1.818787, 
    1.818787, 1.818787,
  1.818734, 1.818736, 1.818735, 1.818737, 1.818736, 1.818737, 1.818734, 
    1.818736, 1.818735, 1.818734, 1.81874, 1.818737, 1.818743, 1.818741, 
    1.818746, 1.818743, 1.818747, 1.818746, 1.818749, 1.818748, 1.818751, 
    1.818749, 1.818753, 1.818751, 1.818751, 1.818749, 1.818738, 1.81874, 
    1.818738, 1.818738, 1.818738, 1.818736, 1.818735, 1.818733, 1.818734, 
    1.818735, 1.818738, 1.818737, 1.818739, 1.818739, 1.818742, 1.818741, 
    1.818745, 1.818744, 1.818748, 1.818747, 1.818748, 1.818748, 1.818748, 
    1.818747, 1.818747, 1.818746, 1.818741, 1.818743, 1.818738, 1.818736, 
    1.818734, 1.818733, 1.818733, 1.818733, 1.818735, 1.818737, 1.818738, 
    1.818739, 1.818739, 1.818742, 1.818743, 1.818746, 1.818745, 1.818746, 
    1.818747, 1.818748, 1.818748, 1.818749, 1.818746, 1.818748, 1.818745, 
    1.818746, 1.81874, 1.818737, 1.818736, 1.818735, 1.818733, 1.818735, 
    1.818734, 1.818735, 1.818736, 1.818736, 1.818739, 1.818738, 1.818743, 
    1.818741, 1.818747, 1.818745, 1.818747, 1.818746, 1.818748, 1.818746, 
    1.818749, 1.81875, 1.818749, 1.818751, 1.818746, 1.818748, 1.818736, 
    1.818736, 1.818736, 1.818735, 1.818735, 1.818733, 1.818735, 1.818735, 
    1.818736, 1.818737, 1.818738, 1.81874, 1.818741, 1.818744, 1.818745, 
    1.818747, 1.818746, 1.818747, 1.818746, 1.818746, 1.818749, 1.818747, 
    1.81875, 1.81875, 1.818749, 1.81875, 1.818736, 1.818736, 1.818734, 
    1.818735, 1.818733, 1.818734, 1.818735, 1.818738, 1.818738, 1.818739, 
    1.81874, 1.818741, 1.818743, 1.818745, 1.818747, 1.818747, 1.818747, 
    1.818747, 1.818746, 1.818748, 1.818748, 1.818747, 1.81875, 1.818749, 
    1.81875, 1.81875, 1.818736, 1.818736, 1.818736, 1.818737, 1.818736, 
    1.818738, 1.818739, 1.818742, 1.818741, 1.818743, 1.818741, 1.818741, 
    1.818743, 1.818741, 1.818745, 1.818743, 1.818747, 1.818745, 1.818748, 
    1.818747, 1.818748, 1.818749, 1.81875, 1.818751, 1.818751, 1.818752, 
    1.818738, 1.818738, 1.818738, 1.818739, 1.81874, 1.818741, 1.818744, 
    1.818743, 1.818745, 1.818745, 1.818742, 1.818744, 1.818739, 1.81874, 
    1.818739, 1.818738, 1.818743, 1.81874, 1.818745, 1.818744, 1.818748, 
    1.818746, 1.818751, 1.818753, 1.818754, 1.818756, 1.818739, 1.818738, 
    1.818739, 1.818741, 1.818742, 1.818744, 1.818744, 1.818745, 1.818745, 
    1.818746, 1.818745, 1.818746, 1.81874, 1.818743, 1.818738, 1.81874, 
    1.818741, 1.81874, 1.818743, 1.818743, 1.818746, 1.818745, 1.818752, 
    1.818749, 1.818758, 1.818755, 1.818738, 1.818739, 1.818742, 1.81874, 
    1.818744, 1.818745, 1.818746, 1.818747, 1.818747, 1.818748, 1.818747, 
    1.818748, 1.818744, 1.818746, 1.818741, 1.818742, 1.818742, 1.818741, 
    1.818743, 1.818745, 1.818745, 1.818745, 1.818747, 1.818744, 1.818753, 
    1.818747, 1.81874, 1.818741, 1.818742, 1.818741, 1.818745, 1.818744, 
    1.818748, 1.818747, 1.818748, 1.818747, 1.818747, 1.818746, 1.818745, 
    1.818744, 1.818742, 1.818741, 1.818741, 1.818743, 1.818745, 1.818747, 
    1.818747, 1.818748, 1.818744, 1.818746, 1.818745, 1.818747, 1.818743, 
    1.818746, 1.818742, 1.818742, 1.818744, 1.818746, 1.818746, 1.818747, 
    1.818747, 1.818745, 1.818745, 1.818743, 1.818743, 1.818742, 1.818742, 
    1.818742, 1.818743, 1.818745, 1.818747, 1.818749, 1.818749, 1.818751, 
    1.81875, 1.818753, 1.81875, 1.818754, 1.818746, 1.81875, 1.818744, 
    1.818744, 1.818745, 1.818748, 1.818747, 1.818749, 1.818745, 1.818743, 
    1.818742, 1.818741, 1.818742, 1.818742, 1.818743, 1.818743, 1.818745, 
    1.818744, 1.818747, 1.818749, 1.818752, 1.818754, 1.818757, 1.818758, 
    1.818758, 1.818758,
  1.818684, 1.818686, 1.818685, 1.818687, 1.818686, 1.818687, 1.818684, 
    1.818686, 1.818685, 1.818684, 1.818691, 1.818687, 1.818694, 1.818692, 
    1.818697, 1.818694, 1.818698, 1.818697, 1.8187, 1.818699, 1.818702, 
    1.8187, 1.818704, 1.818702, 1.818702, 1.8187, 1.818688, 1.81869, 
    1.818688, 1.818688, 1.818688, 1.818686, 1.818685, 1.818683, 1.818684, 
    1.818685, 1.818688, 1.818687, 1.81869, 1.81869, 1.818693, 1.818691, 
    1.818696, 1.818695, 1.818699, 1.818698, 1.818699, 1.818699, 1.818699, 
    1.818697, 1.818698, 1.818697, 1.818692, 1.818693, 1.818689, 1.818686, 
    1.818684, 1.818683, 1.818683, 1.818683, 1.818685, 1.818687, 1.818688, 
    1.818689, 1.81869, 1.818692, 1.818694, 1.818697, 1.818696, 1.818697, 
    1.818698, 1.818699, 1.818699, 1.8187, 1.818697, 1.818699, 1.818696, 
    1.818697, 1.81869, 1.818687, 1.818686, 1.818685, 1.818683, 1.818685, 
    1.818684, 1.818686, 1.818686, 1.818686, 1.818689, 1.818688, 1.818694, 
    1.818691, 1.818698, 1.818696, 1.818698, 1.818697, 1.818699, 1.818697, 
    1.8187, 1.818701, 1.8187, 1.818702, 1.818697, 1.818699, 1.818686, 
    1.818686, 1.818686, 1.818685, 1.818685, 1.818683, 1.818685, 1.818685, 
    1.818687, 1.818687, 1.818688, 1.81869, 1.818692, 1.818694, 1.818696, 
    1.818698, 1.818697, 1.818697, 1.818697, 1.818696, 1.8187, 1.818698, 
    1.818702, 1.818701, 1.8187, 1.818701, 1.818686, 1.818686, 1.818684, 
    1.818685, 1.818683, 1.818684, 1.818685, 1.818688, 1.818688, 1.818689, 
    1.81869, 1.818691, 1.818694, 1.818696, 1.818698, 1.818698, 1.818698, 
    1.818698, 1.818697, 1.818698, 1.818699, 1.818698, 1.818701, 1.8187, 
    1.818701, 1.818701, 1.818686, 1.818687, 1.818686, 1.818687, 1.818686, 
    1.818689, 1.818689, 1.818693, 1.818691, 1.818694, 1.818692, 1.818692, 
    1.818694, 1.818692, 1.818696, 1.818693, 1.818698, 1.818695, 1.818698, 
    1.818698, 1.818699, 1.8187, 1.818701, 1.818702, 1.818702, 1.818704, 
    1.818688, 1.818689, 1.818689, 1.81869, 1.81869, 1.818692, 1.818694, 
    1.818694, 1.818695, 1.818696, 1.818693, 1.818695, 1.818689, 1.81869, 
    1.81869, 1.818688, 1.818694, 1.818691, 1.818696, 1.818695, 1.818699, 
    1.818697, 1.818702, 1.818704, 1.818706, 1.818708, 1.818689, 1.818689, 
    1.81869, 1.818691, 1.818693, 1.818695, 1.818695, 1.818695, 1.818696, 
    1.818697, 1.818695, 1.818697, 1.81869, 1.818694, 1.818688, 1.81869, 
    1.818691, 1.818691, 1.818693, 1.818694, 1.818697, 1.818695, 1.818703, 
    1.8187, 1.818709, 1.818707, 1.818688, 1.818689, 1.818692, 1.818691, 
    1.818695, 1.818696, 1.818697, 1.818698, 1.818698, 1.818699, 1.818697, 
    1.818699, 1.818695, 1.818696, 1.818692, 1.818693, 1.818692, 1.818692, 
    1.818694, 1.818695, 1.818696, 1.818696, 1.818698, 1.818695, 1.818704, 
    1.818698, 1.81869, 1.818692, 1.818692, 1.818691, 1.818696, 1.818694, 
    1.818699, 1.818697, 1.818699, 1.818698, 1.818698, 1.818697, 1.818696, 
    1.818694, 1.818693, 1.818691, 1.818692, 1.818693, 1.818696, 1.818698, 
    1.818697, 1.818699, 1.818695, 1.818696, 1.818696, 1.818698, 1.818694, 
    1.818697, 1.818693, 1.818693, 1.818694, 1.818697, 1.818697, 1.818698, 
    1.818697, 1.818696, 1.818695, 1.818694, 1.818694, 1.818693, 1.818692, 
    1.818693, 1.818694, 1.818696, 1.818698, 1.8187, 1.8187, 1.818702, 
    1.818701, 1.818704, 1.818701, 1.818706, 1.818697, 1.818701, 1.818694, 
    1.818695, 1.818696, 1.818699, 1.818698, 1.8187, 1.818695, 1.818693, 
    1.818693, 1.818692, 1.818693, 1.818693, 1.818694, 1.818693, 1.818696, 
    1.818694, 1.818698, 1.818699, 1.818703, 1.818706, 1.818708, 1.818709, 
    1.81871, 1.81871,
  1.818644, 1.818646, 1.818645, 1.818647, 1.818646, 1.818647, 1.818644, 
    1.818646, 1.818645, 1.818644, 1.818651, 1.818647, 1.818654, 1.818652, 
    1.818657, 1.818654, 1.818658, 1.818657, 1.81866, 1.818659, 1.818662, 
    1.81866, 1.818664, 1.818662, 1.818662, 1.81866, 1.818648, 1.81865, 
    1.818648, 1.818648, 1.818648, 1.818646, 1.818645, 1.818643, 1.818644, 
    1.818645, 1.818648, 1.818647, 1.81865, 1.81865, 1.818653, 1.818651, 
    1.818656, 1.818655, 1.818659, 1.818658, 1.818659, 1.818659, 1.818659, 
    1.818657, 1.818658, 1.818657, 1.818652, 1.818653, 1.818649, 1.818646, 
    1.818644, 1.818643, 1.818643, 1.818643, 1.818645, 1.818647, 1.818648, 
    1.818649, 1.81865, 1.818652, 1.818654, 1.818657, 1.818656, 1.818657, 
    1.818658, 1.818659, 1.818659, 1.81866, 1.818657, 1.818659, 1.818656, 
    1.818657, 1.81865, 1.818648, 1.818646, 1.818645, 1.818643, 1.818645, 
    1.818644, 1.818646, 1.818647, 1.818646, 1.818649, 1.818648, 1.818654, 
    1.818651, 1.818658, 1.818656, 1.818658, 1.818657, 1.818659, 1.818657, 
    1.81866, 1.81866, 1.81866, 1.818662, 1.818657, 1.818659, 1.818646, 
    1.818646, 1.818647, 1.818645, 1.818645, 1.818643, 1.818645, 1.818645, 
    1.818647, 1.818647, 1.818648, 1.81865, 1.818652, 1.818654, 1.818656, 
    1.818658, 1.818657, 1.818657, 1.818657, 1.818656, 1.81866, 1.818658, 
    1.818661, 1.818661, 1.81866, 1.818661, 1.818646, 1.818646, 1.818644, 
    1.818645, 1.818643, 1.818645, 1.818645, 1.818648, 1.818648, 1.818649, 
    1.81865, 1.818651, 1.818654, 1.818656, 1.818658, 1.818658, 1.818658, 
    1.818658, 1.818657, 1.818658, 1.818659, 1.818658, 1.818661, 1.81866, 
    1.818661, 1.818661, 1.818646, 1.818647, 1.818646, 1.818647, 1.818646, 
    1.818649, 1.81865, 1.818653, 1.818651, 1.818654, 1.818652, 1.818652, 
    1.818654, 1.818652, 1.818656, 1.818653, 1.818658, 1.818655, 1.818658, 
    1.818658, 1.818659, 1.81866, 1.81866, 1.818662, 1.818662, 1.818663, 
    1.818648, 1.818649, 1.818649, 1.81865, 1.81865, 1.818652, 1.818654, 
    1.818653, 1.818655, 1.818656, 1.818653, 1.818655, 1.818649, 1.81865, 
    1.81865, 1.818648, 1.818654, 1.818651, 1.818656, 1.818655, 1.818659, 
    1.818657, 1.818662, 1.818664, 1.818666, 1.818668, 1.818649, 1.818649, 
    1.81865, 1.818651, 1.818653, 1.818655, 1.818655, 1.818655, 1.818656, 
    1.818657, 1.818655, 1.818657, 1.81865, 1.818654, 1.818648, 1.81865, 
    1.818651, 1.818651, 1.818653, 1.818654, 1.818657, 1.818655, 1.818663, 
    1.81866, 1.818669, 1.818667, 1.818648, 1.818649, 1.818652, 1.818651, 
    1.818655, 1.818656, 1.818657, 1.818658, 1.818658, 1.818658, 1.818657, 
    1.818658, 1.818655, 1.818656, 1.818652, 1.818653, 1.818653, 1.818652, 
    1.818654, 1.818655, 1.818655, 1.818656, 1.818658, 1.818655, 1.818664, 
    1.818658, 1.81865, 1.818652, 1.818652, 1.818651, 1.818656, 1.818654, 
    1.818658, 1.818657, 1.818659, 1.818658, 1.818658, 1.818657, 1.818656, 
    1.818654, 1.818653, 1.818651, 1.818652, 1.818653, 1.818656, 1.818658, 
    1.818657, 1.818659, 1.818655, 1.818656, 1.818656, 1.818658, 1.818653, 
    1.818657, 1.818653, 1.818653, 1.818654, 1.818657, 1.818657, 1.818658, 
    1.818657, 1.818656, 1.818655, 1.818654, 1.818654, 1.818653, 1.818652, 
    1.818653, 1.818654, 1.818656, 1.818658, 1.81866, 1.81866, 1.818662, 
    1.81866, 1.818664, 1.818661, 1.818666, 1.818657, 1.818661, 1.818654, 
    1.818655, 1.818656, 1.818659, 1.818658, 1.81866, 1.818655, 1.818653, 
    1.818653, 1.818652, 1.818653, 1.818653, 1.818654, 1.818653, 1.818656, 
    1.818654, 1.818658, 1.818659, 1.818663, 1.818666, 1.818668, 1.818669, 
    1.818669, 1.81867,
  1.818579, 1.818581, 1.818581, 1.818582, 1.818581, 1.818582, 1.81858, 
    1.818581, 1.81858, 1.818579, 1.818585, 1.818582, 1.818588, 1.818586, 
    1.818591, 1.818588, 1.818591, 1.818591, 1.818593, 1.818592, 1.818595, 
    1.818593, 1.818596, 1.818594, 1.818595, 1.818593, 1.818583, 1.818585, 
    1.818583, 1.818583, 1.818583, 1.818581, 1.818581, 1.818579, 1.818579, 
    1.818581, 1.818583, 1.818582, 1.818584, 1.818584, 1.818587, 1.818586, 
    1.81859, 1.818589, 1.818592, 1.818591, 1.818592, 1.818592, 1.818592, 
    1.818591, 1.818591, 1.81859, 1.818586, 1.818587, 1.818583, 1.818581, 
    1.81858, 1.818579, 1.818579, 1.818579, 1.818581, 1.818582, 1.818583, 
    1.818584, 1.818584, 1.818586, 1.818588, 1.81859, 1.81859, 1.818591, 
    1.818591, 1.818592, 1.818592, 1.818593, 1.81859, 1.818592, 1.818589, 
    1.81859, 1.818585, 1.818582, 1.818582, 1.818581, 1.818579, 1.81858, 
    1.81858, 1.818581, 1.818582, 1.818581, 1.818584, 1.818583, 1.818588, 
    1.818586, 1.818591, 1.81859, 1.818591, 1.818591, 1.818592, 1.818591, 
    1.818593, 1.818594, 1.818593, 1.818594, 1.818591, 1.818592, 1.818581, 
    1.818581, 1.818582, 1.81858, 1.81858, 1.818579, 1.81858, 1.818581, 
    1.818582, 1.818582, 1.818583, 1.818584, 1.818586, 1.818588, 1.81859, 
    1.818591, 1.81859, 1.818591, 1.81859, 1.81859, 1.818593, 1.818591, 
    1.818594, 1.818594, 1.818593, 1.818594, 1.818581, 1.818581, 1.81858, 
    1.818581, 1.818579, 1.81858, 1.818581, 1.818583, 1.818583, 1.818584, 
    1.818585, 1.818586, 1.818588, 1.81859, 1.818591, 1.818591, 1.818591, 
    1.818592, 1.818591, 1.818592, 1.818592, 1.818591, 1.818594, 1.818593, 
    1.818594, 1.818594, 1.818581, 1.818582, 1.818581, 1.818582, 1.818582, 
    1.818584, 1.818584, 1.818587, 1.818586, 1.818588, 1.818586, 1.818586, 
    1.818588, 1.818586, 1.81859, 1.818587, 1.818592, 1.818589, 1.818592, 
    1.818591, 1.818592, 1.818593, 1.818594, 1.818595, 1.818595, 1.818596, 
    1.818583, 1.818583, 1.818583, 1.818584, 1.818585, 1.818586, 1.818588, 
    1.818588, 1.818589, 1.818589, 1.818587, 1.818588, 1.818584, 1.818585, 
    1.818584, 1.818583, 1.818588, 1.818585, 1.81859, 1.818588, 1.818593, 
    1.818591, 1.818595, 1.818596, 1.818598, 1.8186, 1.818584, 1.818583, 
    1.818584, 1.818586, 1.818587, 1.818589, 1.818589, 1.818589, 1.81859, 
    1.818591, 1.818589, 1.818591, 1.818585, 1.818588, 1.818583, 1.818585, 
    1.818586, 1.818585, 1.818587, 1.818588, 1.81859, 1.818589, 1.818596, 
    1.818593, 1.818601, 1.818599, 1.818583, 1.818584, 1.818586, 1.818585, 
    1.818589, 1.81859, 1.81859, 1.818591, 1.818591, 1.818592, 1.818591, 
    1.818592, 1.818589, 1.81859, 1.818586, 1.818587, 1.818587, 1.818586, 
    1.818588, 1.818589, 1.818589, 1.81859, 1.818591, 1.818589, 1.818596, 
    1.818592, 1.818585, 1.818586, 1.818586, 1.818586, 1.818589, 1.818588, 
    1.818592, 1.818591, 1.818592, 1.818592, 1.818591, 1.81859, 1.81859, 
    1.818588, 1.818587, 1.818586, 1.818586, 1.818587, 1.818589, 1.818591, 
    1.818591, 1.818592, 1.818588, 1.81859, 1.818589, 1.818591, 1.818588, 
    1.818591, 1.818587, 1.818587, 1.818588, 1.81859, 1.818591, 1.818591, 
    1.818591, 1.818589, 1.818589, 1.818588, 1.818588, 1.818587, 1.818586, 
    1.818587, 1.818588, 1.818589, 1.818591, 1.818593, 1.818593, 1.818595, 
    1.818594, 1.818596, 1.818594, 1.818598, 1.818591, 1.818594, 1.818588, 
    1.818589, 1.81859, 1.818592, 1.818591, 1.818593, 1.818589, 1.818587, 
    1.818587, 1.818586, 1.818587, 1.818587, 1.818588, 1.818587, 1.818589, 
    1.818588, 1.818591, 1.818593, 1.818596, 1.818598, 1.8186, 1.818601, 
    1.818601, 1.818601,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2_HR_S1 =
  1.327509e-09, 1.333351e-09, 1.332215e-09, 1.336927e-09, 1.334313e-09, 
    1.337398e-09, 1.328693e-09, 1.333583e-09, 1.330462e-09, 1.328035e-09, 
    1.346071e-09, 1.337137e-09, 1.35535e-09, 1.349652e-09, 1.363964e-09, 
    1.354463e-09, 1.36588e-09, 1.36369e-09, 1.370281e-09, 1.368393e-09, 
    1.376823e-09, 1.371152e-09, 1.381193e-09, 1.375469e-09, 1.376364e-09, 
    1.370965e-09, 1.338935e-09, 1.344959e-09, 1.338578e-09, 1.339437e-09, 
    1.339051e-09, 1.334367e-09, 1.332007e-09, 1.327063e-09, 1.32796e-09, 
    1.331591e-09, 1.339823e-09, 1.337029e-09, 1.344071e-09, 1.343912e-09, 
    1.351752e-09, 1.348217e-09, 1.361394e-09, 1.357649e-09, 1.368472e-09, 
    1.36575e-09, 1.368344e-09, 1.367557e-09, 1.368354e-09, 1.364362e-09, 
    1.366073e-09, 1.36256e-09, 1.348879e-09, 1.3529e-09, 1.340908e-09, 
    1.333698e-09, 1.328908e-09, 1.325509e-09, 1.32599e-09, 1.326906e-09, 
    1.331613e-09, 1.336038e-09, 1.33941e-09, 1.341666e-09, 1.343889e-09, 
    1.350618e-09, 1.354178e-09, 1.362152e-09, 1.360713e-09, 1.36315e-09, 
    1.365479e-09, 1.369389e-09, 1.368745e-09, 1.370468e-09, 1.363086e-09, 
    1.367992e-09, 1.359893e-09, 1.362108e-09, 1.344494e-09, 1.337783e-09, 
    1.33493e-09, 1.332433e-09, 1.326359e-09, 1.330554e-09, 1.3289e-09, 
    1.332834e-09, 1.335334e-09, 1.334098e-09, 1.341728e-09, 1.338762e-09, 
    1.354389e-09, 1.347658e-09, 1.365208e-09, 1.361008e-09, 1.366214e-09, 
    1.363557e-09, 1.368109e-09, 1.364013e-09, 1.371109e-09, 1.372654e-09, 
    1.371598e-09, 1.375655e-09, 1.363786e-09, 1.368344e-09, 1.334063e-09, 
    1.334265e-09, 1.335204e-09, 1.331075e-09, 1.330822e-09, 1.327038e-09, 
    1.330405e-09, 1.331839e-09, 1.335479e-09, 1.337632e-09, 1.339679e-09, 
    1.344179e-09, 1.349204e-09, 1.356232e-09, 1.36128e-09, 1.364664e-09, 
    1.362589e-09, 1.364421e-09, 1.362373e-09, 1.361413e-09, 1.372075e-09, 
    1.366089e-09, 1.375071e-09, 1.374574e-09, 1.370509e-09, 1.37463e-09, 
    1.334406e-09, 1.333246e-09, 1.329217e-09, 1.33237e-09, 1.326626e-09, 
    1.329841e-09, 1.33169e-09, 1.338824e-09, 1.340391e-09, 1.341844e-09, 
    1.344714e-09, 1.348398e-09, 1.35486e-09, 1.360482e-09, 1.365615e-09, 
    1.365238e-09, 1.365371e-09, 1.366517e-09, 1.363677e-09, 1.366984e-09, 
    1.367539e-09, 1.366088e-09, 1.374508e-09, 1.372102e-09, 1.374563e-09, 
    1.372997e-09, 1.333623e-09, 1.335576e-09, 1.334521e-09, 1.336505e-09, 
    1.335107e-09, 1.341322e-09, 1.343185e-09, 1.351904e-09, 1.348326e-09, 
    1.35402e-09, 1.348904e-09, 1.349811e-09, 1.354206e-09, 1.34918e-09, 
    1.360172e-09, 1.35272e-09, 1.366562e-09, 1.359121e-09, 1.367028e-09, 
    1.365592e-09, 1.36797e-09, 1.370099e-09, 1.372778e-09, 1.377721e-09, 
    1.376576e-09, 1.38071e-09, 1.338486e-09, 1.341019e-09, 1.340796e-09, 
    1.343446e-09, 1.345406e-09, 1.349654e-09, 1.356467e-09, 1.353905e-09, 
    1.358608e-09, 1.359553e-09, 1.352407e-09, 1.356794e-09, 1.342713e-09, 
    1.344989e-09, 1.343634e-09, 1.338686e-09, 1.354495e-09, 1.346382e-09, 
    1.361364e-09, 1.356969e-09, 1.369796e-09, 1.363417e-09, 1.375946e-09, 
    1.381303e-09, 1.386344e-09, 1.392235e-09, 1.342401e-09, 1.34068e-09, 
    1.343761e-09, 1.348024e-09, 1.351979e-09, 1.357237e-09, 1.357775e-09, 
    1.35876e-09, 1.361311e-09, 1.363456e-09, 1.359071e-09, 1.363994e-09, 
    1.345516e-09, 1.3552e-09, 1.34003e-09, 1.344598e-09, 1.347772e-09, 
    1.34638e-09, 1.353612e-09, 1.355317e-09, 1.362244e-09, 1.358663e-09, 
    1.379981e-09, 1.370549e-09, 1.396721e-09, 1.389407e-09, 1.340079e-09, 
    1.342395e-09, 1.350455e-09, 1.34662e-09, 1.357588e-09, 1.360287e-09, 
    1.362482e-09, 1.365287e-09, 1.36559e-09, 1.367252e-09, 1.364528e-09, 
    1.367145e-09, 1.357248e-09, 1.36167e-09, 1.349534e-09, 1.352488e-09, 
    1.351129e-09, 1.349638e-09, 1.354239e-09, 1.35914e-09, 1.359245e-09, 
    1.360816e-09, 1.365246e-09, 1.357632e-09, 1.381199e-09, 1.366645e-09, 
    1.34492e-09, 1.349381e-09, 1.350018e-09, 1.34829e-09, 1.360017e-09, 
    1.355768e-09, 1.367212e-09, 1.364119e-09, 1.369186e-09, 1.366668e-09, 
    1.366298e-09, 1.363063e-09, 1.36105e-09, 1.355963e-09, 1.351823e-09, 
    1.348541e-09, 1.349304e-09, 1.35291e-09, 1.35944e-09, 1.365618e-09, 
    1.364264e-09, 1.368801e-09, 1.356792e-09, 1.361828e-09, 1.359882e-09, 
    1.364956e-09, 1.353837e-09, 1.363306e-09, 1.351416e-09, 1.352459e-09, 
    1.355683e-09, 1.36217e-09, 1.363604e-09, 1.365137e-09, 1.364191e-09, 
    1.359606e-09, 1.358854e-09, 1.355605e-09, 1.354708e-09, 1.352232e-09, 
    1.350182e-09, 1.352055e-09, 1.354022e-09, 1.359608e-09, 1.364641e-09, 
    1.37013e-09, 1.371473e-09, 1.377885e-09, 1.372665e-09, 1.38128e-09, 
    1.373956e-09, 1.386633e-09, 1.363855e-09, 1.373741e-09, 1.35583e-09, 
    1.35776e-09, 1.36125e-09, 1.369254e-09, 1.364933e-09, 1.369987e-09, 
    1.358825e-09, 1.353034e-09, 1.351536e-09, 1.34874e-09, 1.3516e-09, 
    1.351367e-09, 1.354103e-09, 1.353224e-09, 1.359793e-09, 1.356264e-09, 
    1.366289e-09, 1.369947e-09, 1.380277e-09, 1.38661e-09, 1.393056e-09, 
    1.395902e-09, 1.396768e-09, 1.39713e-09 ;

 SOIL2_HR_S3 =
  9.482209e-11, 9.523934e-11, 9.515823e-11, 9.549478e-11, 9.530808e-11, 
    9.552846e-11, 9.490668e-11, 9.525591e-11, 9.503297e-11, 9.485965e-11, 
    9.614792e-11, 9.550979e-11, 9.68107e-11, 9.640374e-11, 9.742602e-11, 
    9.674738e-11, 9.756286e-11, 9.740643e-11, 9.787721e-11, 9.774234e-11, 
    9.834452e-11, 9.793946e-11, 9.865665e-11, 9.824778e-11, 9.831175e-11, 
    9.79261e-11, 9.56382e-11, 9.606847e-11, 9.561271e-11, 9.567407e-11, 
    9.564653e-11, 9.531195e-11, 9.514334e-11, 9.479019e-11, 9.48543e-11, 
    9.511367e-11, 9.570165e-11, 9.550206e-11, 9.600507e-11, 9.599371e-11, 
    9.655372e-11, 9.630122e-11, 9.724245e-11, 9.697494e-11, 9.774797e-11, 
    9.755356e-11, 9.773884e-11, 9.768265e-11, 9.773957e-11, 9.745445e-11, 
    9.757661e-11, 9.732572e-11, 9.634851e-11, 9.663571e-11, 9.577915e-11, 
    9.526412e-11, 9.4922e-11, 9.467923e-11, 9.471356e-11, 9.477898e-11, 
    9.511519e-11, 9.543129e-11, 9.567217e-11, 9.583331e-11, 9.599208e-11, 
    9.647268e-11, 9.672703e-11, 9.729655e-11, 9.719376e-11, 9.736788e-11, 
    9.753422e-11, 9.781349e-11, 9.776752e-11, 9.789057e-11, 9.736328e-11, 
    9.771373e-11, 9.713522e-11, 9.729344e-11, 9.603528e-11, 9.55559e-11, 
    9.535218e-11, 9.517382e-11, 9.473994e-11, 9.503957e-11, 9.492146e-11, 
    9.520246e-11, 9.538101e-11, 9.52927e-11, 9.583772e-11, 9.562583e-11, 
    9.674211e-11, 9.626129e-11, 9.751482e-11, 9.721485e-11, 9.758672e-11, 
    9.739697e-11, 9.772209e-11, 9.742948e-11, 9.793636e-11, 9.804674e-11, 
    9.797131e-11, 9.826104e-11, 9.741326e-11, 9.773884e-11, 9.529023e-11, 
    9.530463e-11, 9.537172e-11, 9.507678e-11, 9.505874e-11, 9.478843e-11, 
    9.502894e-11, 9.513137e-11, 9.539135e-11, 9.554515e-11, 9.569134e-11, 
    9.601276e-11, 9.637174e-11, 9.68737e-11, 9.72343e-11, 9.747603e-11, 
    9.73278e-11, 9.745867e-11, 9.731237e-11, 9.724381e-11, 9.800538e-11, 
    9.757775e-11, 9.821936e-11, 9.818386e-11, 9.78935e-11, 9.818786e-11, 
    9.531474e-11, 9.523186e-11, 9.49441e-11, 9.51693e-11, 9.475899e-11, 
    9.498867e-11, 9.512073e-11, 9.563027e-11, 9.574221e-11, 9.584602e-11, 
    9.605104e-11, 9.631415e-11, 9.677571e-11, 9.71773e-11, 9.75439e-11, 
    9.751704e-11, 9.752649e-11, 9.760839e-11, 9.740553e-11, 9.764169e-11, 
    9.768134e-11, 9.75777e-11, 9.81791e-11, 9.800729e-11, 9.818311e-11, 
    9.807123e-11, 9.52588e-11, 9.539826e-11, 9.53229e-11, 9.546461e-11, 
    9.536478e-11, 9.58087e-11, 9.59418e-11, 9.656457e-11, 9.630897e-11, 
    9.671574e-11, 9.635029e-11, 9.641504e-11, 9.672903e-11, 9.637004e-11, 
    9.715517e-11, 9.662289e-11, 9.761157e-11, 9.708006e-11, 9.764489e-11, 
    9.754231e-11, 9.771213e-11, 9.786423e-11, 9.805558e-11, 9.840864e-11, 
    9.832688e-11, 9.862215e-11, 9.560616e-11, 9.578705e-11, 9.577112e-11, 
    9.596042e-11, 9.610041e-11, 9.640384e-11, 9.68905e-11, 9.670749e-11, 
    9.704346e-11, 9.71109e-11, 9.660048e-11, 9.691389e-11, 9.590811e-11, 
    9.607062e-11, 9.597385e-11, 9.562044e-11, 9.674968e-11, 9.617016e-11, 
    9.724026e-11, 9.692632e-11, 9.784255e-11, 9.73869e-11, 9.828188e-11, 
    9.866449e-11, 9.902455e-11, 9.944538e-11, 9.588577e-11, 9.576286e-11, 
    9.598293e-11, 9.628742e-11, 9.65699e-11, 9.694547e-11, 9.698389e-11, 
    9.705426e-11, 9.72365e-11, 9.738974e-11, 9.707651e-11, 9.742814e-11, 
    9.610832e-11, 9.679997e-11, 9.571639e-11, 9.60427e-11, 9.626946e-11, 
    9.616998e-11, 9.668658e-11, 9.680833e-11, 9.730311e-11, 9.704734e-11, 
    9.857007e-11, 9.789637e-11, 9.976577e-11, 9.924336e-11, 9.571992e-11, 
    9.588534e-11, 9.646108e-11, 9.618715e-11, 9.697054e-11, 9.716337e-11, 
    9.732012e-11, 9.752051e-11, 9.754214e-11, 9.766087e-11, 9.746631e-11, 
    9.765318e-11, 9.694628e-11, 9.726218e-11, 9.639527e-11, 9.660627e-11, 
    9.65092e-11, 9.640273e-11, 9.673134e-11, 9.708145e-11, 9.708891e-11, 
    9.720118e-11, 9.751755e-11, 9.697371e-11, 9.865705e-11, 9.761748e-11, 
    9.606573e-11, 9.638438e-11, 9.642988e-11, 9.630644e-11, 9.714404e-11, 
    9.684056e-11, 9.765798e-11, 9.743705e-11, 9.779903e-11, 9.761916e-11, 
    9.75927e-11, 9.736167e-11, 9.721784e-11, 9.685447e-11, 9.655881e-11, 
    9.632434e-11, 9.637886e-11, 9.663641e-11, 9.710286e-11, 9.754411e-11, 
    9.744745e-11, 9.777152e-11, 9.691374e-11, 9.727343e-11, 9.713442e-11, 
    9.749689e-11, 9.670263e-11, 9.737903e-11, 9.652974e-11, 9.66042e-11, 
    9.683453e-11, 9.729784e-11, 9.740032e-11, 9.750976e-11, 9.744223e-11, 
    9.71147e-11, 9.706103e-11, 9.682893e-11, 9.676485e-11, 9.658799e-11, 
    9.644157e-11, 9.657535e-11, 9.671584e-11, 9.711483e-11, 9.747439e-11, 
    9.78664e-11, 9.796233e-11, 9.842039e-11, 9.804753e-11, 9.866283e-11, 
    9.813974e-11, 9.904524e-11, 9.741821e-11, 9.812433e-11, 9.6845e-11, 
    9.698282e-11, 9.723212e-11, 9.780387e-11, 9.749519e-11, 9.785618e-11, 
    9.705893e-11, 9.66453e-11, 9.653827e-11, 9.63386e-11, 9.654284e-11, 
    9.652622e-11, 9.672166e-11, 9.665885e-11, 9.712808e-11, 9.687603e-11, 
    9.759203e-11, 9.785332e-11, 9.85912e-11, 9.904355e-11, 9.950399e-11, 
    9.970727e-11, 9.976914e-11, 9.979501e-11 ;

 SOIL3C =
  5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782611, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782613, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782613, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782613, 5.782613, 
    5.782613, 5.782613 ;

 SOIL3C_TO_SOIL1C =
  2.6178e-11, 2.629317e-11, 2.627078e-11, 2.636367e-11, 2.631214e-11, 
    2.637296e-11, 2.620134e-11, 2.629774e-11, 2.62362e-11, 2.618836e-11, 
    2.654394e-11, 2.636781e-11, 2.672688e-11, 2.661455e-11, 2.689672e-11, 
    2.67094e-11, 2.693448e-11, 2.689131e-11, 2.702125e-11, 2.698402e-11, 
    2.715023e-11, 2.703843e-11, 2.723639e-11, 2.712353e-11, 2.714119e-11, 
    2.703474e-11, 2.640325e-11, 2.652202e-11, 2.639622e-11, 2.641315e-11, 
    2.640555e-11, 2.63132e-11, 2.626667e-11, 2.616919e-11, 2.618689e-11, 
    2.625848e-11, 2.642077e-11, 2.636568e-11, 2.650452e-11, 2.650138e-11, 
    2.665595e-11, 2.658626e-11, 2.684605e-11, 2.677221e-11, 2.698558e-11, 
    2.693192e-11, 2.698306e-11, 2.696755e-11, 2.698326e-11, 2.690456e-11, 
    2.693828e-11, 2.686903e-11, 2.659931e-11, 2.667858e-11, 2.644216e-11, 
    2.63e-11, 2.620557e-11, 2.613857e-11, 2.614804e-11, 2.61661e-11, 
    2.62589e-11, 2.634614e-11, 2.641263e-11, 2.645711e-11, 2.650093e-11, 
    2.663358e-11, 2.670379e-11, 2.686098e-11, 2.683261e-11, 2.688067e-11, 
    2.692658e-11, 2.700366e-11, 2.699098e-11, 2.702494e-11, 2.68794e-11, 
    2.697613e-11, 2.681645e-11, 2.686012e-11, 2.651286e-11, 2.638054e-11, 
    2.632431e-11, 2.627508e-11, 2.615532e-11, 2.623803e-11, 2.620542e-11, 
    2.628298e-11, 2.633227e-11, 2.630789e-11, 2.645833e-11, 2.639984e-11, 
    2.670795e-11, 2.657524e-11, 2.692123e-11, 2.683843e-11, 2.694107e-11, 
    2.68887e-11, 2.697844e-11, 2.689767e-11, 2.703758e-11, 2.706804e-11, 
    2.704722e-11, 2.712719e-11, 2.689319e-11, 2.698306e-11, 2.630721e-11, 
    2.631118e-11, 2.63297e-11, 2.62483e-11, 2.624331e-11, 2.616871e-11, 
    2.623509e-11, 2.626336e-11, 2.633512e-11, 2.637757e-11, 2.641792e-11, 
    2.650664e-11, 2.660572e-11, 2.674427e-11, 2.68438e-11, 2.691052e-11, 
    2.686961e-11, 2.690573e-11, 2.686535e-11, 2.684642e-11, 2.705663e-11, 
    2.69386e-11, 2.711569e-11, 2.710589e-11, 2.702574e-11, 2.710699e-11, 
    2.631398e-11, 2.62911e-11, 2.621167e-11, 2.627383e-11, 2.616058e-11, 
    2.622398e-11, 2.626043e-11, 2.640107e-11, 2.643196e-11, 2.646062e-11, 
    2.65172e-11, 2.658983e-11, 2.671722e-11, 2.682807e-11, 2.692925e-11, 
    2.692184e-11, 2.692445e-11, 2.694705e-11, 2.689106e-11, 2.695624e-11, 
    2.696719e-11, 2.693858e-11, 2.710458e-11, 2.705715e-11, 2.710568e-11, 
    2.70748e-11, 2.629853e-11, 2.633703e-11, 2.631623e-11, 2.635534e-11, 
    2.632779e-11, 2.645032e-11, 2.648705e-11, 2.665894e-11, 2.65884e-11, 
    2.670067e-11, 2.65998e-11, 2.661768e-11, 2.670434e-11, 2.660525e-11, 
    2.682196e-11, 2.667504e-11, 2.694793e-11, 2.680123e-11, 2.695712e-11, 
    2.692881e-11, 2.697569e-11, 2.701767e-11, 2.707048e-11, 2.716793e-11, 
    2.714536e-11, 2.722686e-11, 2.639441e-11, 2.644434e-11, 2.643994e-11, 
    2.649219e-11, 2.653083e-11, 2.661458e-11, 2.674891e-11, 2.669839e-11, 
    2.679112e-11, 2.680974e-11, 2.666886e-11, 2.675536e-11, 2.647775e-11, 
    2.652261e-11, 2.64959e-11, 2.639835e-11, 2.671004e-11, 2.655008e-11, 
    2.684544e-11, 2.675879e-11, 2.701168e-11, 2.688592e-11, 2.713294e-11, 
    2.723855e-11, 2.733793e-11, 2.745408e-11, 2.647159e-11, 2.643766e-11, 
    2.64984e-11, 2.658245e-11, 2.666042e-11, 2.676408e-11, 2.677468e-11, 
    2.679411e-11, 2.684441e-11, 2.68867e-11, 2.680025e-11, 2.68973e-11, 
    2.653302e-11, 2.672392e-11, 2.642484e-11, 2.65149e-11, 2.657749e-11, 
    2.655003e-11, 2.669262e-11, 2.672623e-11, 2.686279e-11, 2.67922e-11, 
    2.721249e-11, 2.702654e-11, 2.754251e-11, 2.739832e-11, 2.642581e-11, 
    2.647147e-11, 2.663038e-11, 2.655477e-11, 2.6771e-11, 2.682422e-11, 
    2.686749e-11, 2.69228e-11, 2.692877e-11, 2.696154e-11, 2.690784e-11, 
    2.695942e-11, 2.67643e-11, 2.685149e-11, 2.661222e-11, 2.667046e-11, 
    2.664366e-11, 2.661428e-11, 2.670498e-11, 2.680161e-11, 2.680367e-11, 
    2.683466e-11, 2.692198e-11, 2.677187e-11, 2.723649e-11, 2.694956e-11, 
    2.652126e-11, 2.660921e-11, 2.662177e-11, 2.65877e-11, 2.681889e-11, 
    2.673512e-11, 2.696074e-11, 2.689976e-11, 2.699967e-11, 2.695002e-11, 
    2.694272e-11, 2.687896e-11, 2.683926e-11, 2.673896e-11, 2.665736e-11, 
    2.659264e-11, 2.660769e-11, 2.667878e-11, 2.680752e-11, 2.692931e-11, 
    2.690263e-11, 2.699208e-11, 2.675532e-11, 2.68546e-11, 2.681623e-11, 
    2.691628e-11, 2.669705e-11, 2.688375e-11, 2.664933e-11, 2.666989e-11, 
    2.673346e-11, 2.686134e-11, 2.688962e-11, 2.691983e-11, 2.690119e-11, 
    2.681079e-11, 2.679598e-11, 2.673191e-11, 2.671423e-11, 2.666541e-11, 
    2.6625e-11, 2.666192e-11, 2.67007e-11, 2.681082e-11, 2.691007e-11, 
    2.701827e-11, 2.704474e-11, 2.717117e-11, 2.706826e-11, 2.723809e-11, 
    2.709371e-11, 2.734364e-11, 2.689456e-11, 2.708946e-11, 2.673635e-11, 
    2.677439e-11, 2.68432e-11, 2.700101e-11, 2.691581e-11, 2.701545e-11, 
    2.679539e-11, 2.668123e-11, 2.665169e-11, 2.659658e-11, 2.665295e-11, 
    2.664836e-11, 2.67023e-11, 2.668497e-11, 2.681448e-11, 2.674491e-11, 
    2.694254e-11, 2.701466e-11, 2.721832e-11, 2.734317e-11, 2.747026e-11, 
    2.752636e-11, 2.754344e-11, 2.755058e-11 ;

 SOIL3C_vr =
  20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009,
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00007, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00007, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00007, 20.00008, 20.00007, 20.00008, 20.00007, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N =
  0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692 ;

 SOIL3N_TNDNCY_VERT_TRANS =
  -2.569961e-21, -7.709882e-21, 5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -7.709882e-21, -5.139921e-21, -7.709882e-21, 1.027984e-20, -5.139921e-21, 
    -7.709882e-21, -2.569961e-21, -1.541976e-20, -2.569961e-21, 
    -2.569961e-21, -5.139921e-21, -1.28498e-20, 1.541976e-20, -1.027984e-20, 
    1.541976e-20, -5.139921e-21, -5.139921e-21, 1.003089e-36, 1.027984e-20, 
    1.027984e-20, -1.003089e-36, -2.569961e-21, -5.139921e-21, -1.798972e-20, 
    5.139921e-21, -2.569961e-21, -1.027984e-20, 2.569961e-21, -2.569961e-21, 
    -1.027984e-20, -1.027984e-20, -1.798972e-20, 1.28498e-20, -1.027984e-20, 
    -1.003089e-36, -1.541976e-20, -7.709882e-21, -2.569961e-21, 
    -2.569961e-21, 1.027984e-20, 0, -5.139921e-21, 0, 2.569961e-21, 
    7.709882e-21, 5.139921e-21, 1.003089e-36, 5.139921e-21, -7.709882e-21, 
    7.709882e-21, -1.003089e-36, -5.139921e-21, -1.027984e-20, -2.569961e-21, 
    5.139921e-21, 7.709882e-21, 0, 1.027984e-20, 2.569961e-21, 0, 
    1.027984e-20, -2.569961e-21, 7.709882e-21, 1.28498e-20, 0, 2.569961e-21, 
    -1.003089e-36, 1.541976e-20, 2.569961e-21, -5.139921e-21, -7.709882e-21, 
    7.709882e-21, 2.569961e-20, -1.28498e-20, -1.541976e-20, 2.569961e-21, 
    1.027984e-20, -1.027984e-20, -7.709882e-21, 1.28498e-20, 7.709882e-21, 0, 
    -7.709882e-21, -1.027984e-20, 7.709882e-21, -2.312965e-20, -1.28498e-20, 
    2.569961e-21, -1.027984e-20, -2.569961e-20, 7.709882e-21, 2.569961e-21, 
    -1.28498e-20, -7.709882e-21, 1.003089e-36, -1.28498e-20, -2.569961e-21, 
    -2.569961e-21, -1.541976e-20, 7.709882e-21, 1.027984e-20, -7.709882e-21, 
    -7.709882e-21, 7.709882e-21, 0, -2.569961e-21, 5.139921e-21, 
    -1.003089e-36, -1.541976e-20, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -1.027984e-20, 2.569961e-21, -1.28498e-20, 7.709882e-21, 
    5.139921e-21, 0, 1.027984e-20, -1.541976e-20, -7.709882e-21, 
    -2.569961e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, -7.709882e-21, 
    2.569961e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, -1.027984e-20, 
    1.003089e-36, -1.541976e-20, 1.027984e-20, 1.003089e-36, -1.027984e-20, 
    -1.027984e-20, 5.139921e-21, -1.541976e-20, 0, -5.139921e-21, 
    1.027984e-20, -2.569961e-21, -5.139921e-21, 1.541976e-20, 0, 
    -2.569961e-21, 2.569961e-21, 2.569961e-21, -1.28498e-20, 2.569961e-21, 
    -5.139921e-21, 1.027984e-20, -2.569961e-21, 1.027984e-20, 1.541976e-20, 
    -7.709882e-21, 1.003089e-36, -5.139921e-21, 7.709882e-21, 1.28498e-20, 
    -1.003089e-36, -1.003089e-36, -1.28498e-20, -2.569961e-21, 2.569961e-21, 
    2.569961e-21, -5.139921e-21, -5.139921e-21, 1.28498e-20, 0, 7.709882e-21, 
    1.027984e-20, -2.569961e-21, 2.569961e-21, 5.139921e-21, -5.139921e-21, 
    2.569961e-21, 1.28498e-20, -5.139921e-21, -2.055969e-20, -1.003089e-36, 
    -2.569961e-21, 0, -1.027984e-20, 1.027984e-20, 1.541976e-20, 
    -5.139921e-21, -2.569961e-21, 1.003089e-36, -7.709882e-21, -5.139921e-21, 
    -2.569961e-21, 1.28498e-20, -5.139921e-21, -2.569961e-21, 1.541976e-20, 
    7.709882e-21, -2.569961e-21, -1.798972e-20, -5.139921e-21, -1.003089e-36, 
    5.139921e-21, 7.709882e-21, 2.569961e-21, 5.139921e-21, 2.569961e-21, 
    1.027984e-20, 7.709882e-21, 2.569961e-21, 1.28498e-20, -2.569961e-21, 
    1.541976e-20, -7.709882e-21, 1.027984e-20, 1.003089e-36, -1.003089e-36, 
    2.569961e-21, -1.027984e-20, 2.569961e-21, 2.312965e-20, -1.541976e-20, 
    1.541976e-20, 0, -1.027984e-20, -1.027984e-20, -1.027984e-20, 
    2.055969e-20, 7.709882e-21, -7.709882e-21, 1.28498e-20, 7.709882e-21, 0, 
    1.28498e-20, -2.569961e-20, -2.569961e-21, 1.027984e-20, -2.569961e-21, 
    1.027984e-20, -1.28498e-20, -2.569961e-21, -2.569961e-21, -1.027984e-20, 
    1.027984e-20, -1.027984e-20, 1.28498e-20, -1.28498e-20, 2.569961e-21, 
    -1.003089e-36, 2.569961e-21, -7.709882e-21, 2.569961e-21, -7.709882e-21, 
    1.003089e-36, 5.139921e-21, -1.003089e-36, -1.027984e-20, 5.139921e-21, 
    -5.139921e-21, 7.709882e-21, 2.826957e-20, 7.709882e-21, -7.709882e-21, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, -7.709882e-21, -1.541976e-20, 
    7.709882e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, 1.027984e-20, 
    -1.541976e-20, 1.541976e-20, 1.003089e-36, 0, 5.139921e-21, 
    -1.003089e-36, 7.709882e-21, -1.027984e-20, 1.541976e-20, 1.027984e-20, 
    2.569961e-21, -1.027984e-20, 1.798972e-20, -7.709882e-21, -7.709882e-21, 
    5.139921e-21, 1.027984e-20, 2.312965e-20, 0, 1.003089e-36, 1.027984e-20, 
    1.541976e-20, 5.139921e-21, -5.139921e-21, -2.569961e-21, 1.798972e-20, 
    -7.709882e-21, 1.28498e-20, 7.709882e-21, 5.139921e-21, 5.139921e-21, 
    -1.027984e-20, -1.027984e-20, 5.139921e-21, 7.709882e-21, 1.003089e-36, 
    1.027984e-20, -7.709882e-21, -2.569961e-21, 1.027984e-20, 1.027984e-20, 
    -1.027984e-20, 1.027984e-20, 1.003089e-36, 7.709882e-21, -1.541976e-20, 
    7.709882e-21, -1.798972e-20, 7.709882e-21, -7.709882e-21, -2.569961e-21, 
    -1.027984e-20, 5.139921e-21, 2.569961e-21, 1.027984e-20, -2.569961e-21, 
    5.139921e-21, 1.798972e-20, 1.28498e-20, -1.28498e-20,
  0, 0, -5.139921e-21, -5.139921e-21, 1.027984e-20, -1.027984e-20, 
    -5.139921e-21, 2.569961e-21, 7.709882e-21, -2.569961e-21, -1.28498e-20, 
    5.139921e-21, 2.569961e-21, 5.139921e-21, 2.569961e-21, 7.709882e-21, 
    2.569961e-21, -2.569961e-21, 7.709882e-21, -7.709882e-21, 5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 2.569961e-21, 2.569961e-21, 7.709882e-21, 
    -2.569961e-21, -7.709882e-21, -7.709882e-21, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 2.569961e-21, -1.541976e-20, 2.569961e-21, -1.027984e-20, 
    2.569961e-21, -5.139921e-21, 1.027984e-20, -7.709882e-21, 1.798972e-20, 
    7.709882e-21, -5.139921e-21, 7.709882e-21, 7.709882e-21, -2.569961e-21, 
    2.569961e-21, -7.709882e-21, 0, -1.027984e-20, -5.139921e-21, 
    1.28498e-20, 0, 0, -5.139921e-21, -1.28498e-20, -5.139921e-21, 
    2.569961e-21, -7.709882e-21, -1.027984e-20, -7.709882e-21, 7.709882e-21, 
    0, 7.709882e-21, 2.569961e-21, 5.139921e-21, 7.709882e-21, -5.139921e-21, 
    -7.709882e-21, -2.569961e-21, 1.027984e-20, 1.027984e-20, 5.139921e-21, 
    -2.569961e-21, 1.027984e-20, -2.569961e-21, 7.709882e-21, -1.027984e-20, 
    5.139921e-21, 5.139921e-21, -2.569961e-21, -2.569961e-21, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, -7.709882e-21, -1.027984e-20, 2.569961e-21, 
    -7.709882e-21, 2.569961e-21, -5.139921e-21, -7.709882e-21, 1.027984e-20, 
    0, -1.28498e-20, 5.139921e-21, -2.569961e-21, 2.569961e-21, 5.139921e-21, 
    7.709882e-21, -5.139921e-21, -1.28498e-20, -7.709882e-21, 0, 
    7.709882e-21, 2.569961e-21, -5.139921e-21, -7.709882e-21, 1.28498e-20, 
    1.027984e-20, 5.139921e-21, 2.569961e-21, 5.139921e-21, 0, 0, 
    -7.709882e-21, -5.139921e-21, 1.027984e-20, 0, -2.569961e-21, 
    1.798972e-20, 5.139921e-21, 1.003089e-36, -5.139921e-21, 2.569961e-21, 
    -7.709882e-21, 1.027984e-20, -1.027984e-20, 1.798972e-20, 7.709882e-21, 
    -7.709882e-21, 1.28498e-20, -5.139921e-21, -2.569961e-21, 2.569961e-21, 
    -7.709882e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, 
    -5.139921e-21, 1.28498e-20, -5.139921e-21, 2.569961e-21, -1.28498e-20, 
    1.541976e-20, -5.139921e-21, -1.027984e-20, 5.139921e-21, -1.28498e-20, 
    7.709882e-21, 5.139921e-21, -7.709882e-21, -1.027984e-20, -5.139921e-21, 
    -1.027984e-20, 0, -1.28498e-20, 1.027984e-20, 1.027984e-20, 
    -7.709882e-21, -1.003089e-36, 5.139921e-21, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 7.709882e-21, 2.569961e-21, 2.569961e-21, -5.139921e-21, 
    0, 2.569961e-21, 1.003089e-36, 0, -1.798972e-20, -5.139921e-21, 
    -5.139921e-21, -1.28498e-20, 2.055969e-20, 7.709882e-21, -5.139921e-21, 
    2.569961e-21, -7.709882e-21, 1.28498e-20, 7.709882e-21, 0, 2.569961e-21, 
    7.709882e-21, -2.569961e-21, 5.139921e-21, 1.28498e-20, 0, 5.139921e-21, 
    7.709882e-21, -2.569961e-21, 0, 1.28498e-20, -7.709882e-21, 0, 
    -1.28498e-20, 7.709882e-21, 1.003089e-36, -2.569961e-21, -7.709882e-21, 
    -2.569961e-21, 2.569961e-21, 7.709882e-21, -1.003089e-36, -1.027984e-20, 
    0, 2.569961e-21, 2.569961e-21, 5.139921e-21, -1.541976e-20, -1.28498e-20, 
    5.139921e-21, -5.139921e-21, 1.28498e-20, -5.139921e-21, 2.569961e-21, 
    -1.027984e-20, 2.569961e-21, -5.139921e-21, 1.027984e-20, 0, 
    5.139921e-21, 2.569961e-21, 1.003089e-36, 2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 1.027984e-20, -1.541976e-20, 2.569961e-21, 2.569961e-21, 
    7.709882e-21, 7.709882e-21, -1.28498e-20, 7.709882e-21, -2.569961e-21, 
    2.569961e-21, -5.139921e-21, 5.139921e-21, 7.709882e-21, 5.139921e-21, 
    -1.027984e-20, -1.003089e-36, -5.139921e-21, 0, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, -1.027984e-20, 1.541976e-20, 7.709882e-21, 
    -2.569961e-21, 2.569961e-21, -1.28498e-20, -2.569961e-21, 2.569961e-21, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, 1.798972e-20, -5.139921e-21, 
    1.003089e-36, 0, -1.541976e-20, 2.569961e-21, -1.027984e-20, 
    -1.541976e-20, -2.569961e-21, -1.027984e-20, 0, 1.027984e-20, 
    -1.28498e-20, 1.28498e-20, -5.139921e-21, 2.569961e-21, 5.139921e-21, 
    5.139921e-21, 1.28498e-20, -7.709882e-21, 5.139921e-21, 1.798972e-20, 
    -2.569961e-21, 0, 2.569961e-21, -5.139921e-21, 5.139921e-21, 
    2.569961e-21, 0, 1.541976e-20, -1.541976e-20, 5.139921e-21, 1.027984e-20, 
    -1.28498e-20, -5.139921e-21, -7.709882e-21, 2.055969e-20, 2.569961e-21, 
    1.541976e-20, -5.139921e-21, -5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -7.709882e-21, 2.569961e-21, 0, -1.003089e-36, 5.139921e-21, 
    7.709882e-21, -5.139921e-21, -5.139921e-21, -5.139921e-21, -5.139921e-21, 
    2.569961e-21, -5.139921e-21, 2.569961e-21, -5.139921e-21, -5.139921e-21, 
    -7.709882e-21, -2.569961e-21, -7.709882e-21, 7.709882e-21, -2.569961e-21, 
    -2.569961e-21, 1.003089e-36, -5.139921e-21, -2.569961e-21, 1.798972e-20, 
    -7.709882e-21, 2.569961e-21, 0, -2.569961e-21, -2.569961e-21, 
    -5.139921e-21, 5.139921e-21,
  -7.709882e-21, -1.28498e-20, 1.027984e-20, 1.003089e-36, -2.569961e-21, 
    -5.139921e-21, 0, -1.798972e-20, 7.709882e-21, 0, -2.569961e-21, 
    -2.569961e-21, 7.709882e-21, 2.569961e-21, 1.798972e-20, -2.055969e-20, 
    -2.569961e-21, 1.027984e-20, -1.003089e-36, -1.027984e-20, 2.569961e-21, 
    2.569961e-21, -1.541976e-20, 5.139921e-21, 5.139921e-21, -7.709882e-21, 
    2.569961e-21, 0, 7.709882e-21, 7.709882e-21, 5.139921e-21, 0, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, 5.139921e-21, 1.28498e-20, 
    1.798972e-20, 1.28498e-20, 1.798972e-20, 0, -2.569961e-21, -1.027984e-20, 
    2.569961e-21, 7.709882e-21, 2.569961e-21, 7.709882e-21, -7.709882e-21, 
    5.139921e-21, -1.541976e-20, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 7.709882e-21, 2.569961e-21, -1.003089e-36, -1.003089e-36, 
    -1.027984e-20, 5.139921e-21, 2.569961e-21, 2.569961e-21, -5.139921e-21, 
    -2.569961e-21, 7.709882e-21, -2.569961e-21, -7.709882e-21, 2.569961e-21, 
    -5.139921e-21, -2.569961e-21, -7.709882e-21, 2.569961e-21, -2.569961e-21, 
    1.28498e-20, -1.003089e-36, 5.139921e-21, -5.139921e-21, 0, 5.139921e-21, 
    -2.569961e-21, -7.709882e-21, 5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -7.709882e-21, -7.709882e-21, 5.139921e-21, -2.569961e-21, 0, 0, 
    1.28498e-20, 1.541976e-20, 7.709882e-21, 0, -7.709882e-21, -2.312965e-20, 
    -5.139921e-21, -2.569961e-21, 1.28498e-20, -2.569961e-21, -1.798972e-20, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, -1.003089e-36, 2.569961e-21, 
    0, 5.139921e-21, -1.003089e-36, 0, 2.569961e-21, -7.709882e-21, 
    2.569961e-21, 2.569961e-21, -1.541976e-20, -2.055969e-20, -7.709882e-21, 
    0, -2.569961e-21, -7.709882e-21, 1.027984e-20, -2.569961e-21, 
    1.003089e-36, 7.709882e-21, 1.28498e-20, -1.003089e-36, -1.027984e-20, 
    7.709882e-21, 2.569961e-21, -5.139921e-21, 2.569961e-21, -5.139921e-21, 
    -1.027984e-20, 1.027984e-20, 7.709882e-21, -5.139921e-21, -7.709882e-21, 
    -1.798972e-20, -5.139921e-21, 1.027984e-20, 7.709882e-21, 1.027984e-20, 
    -2.569961e-21, -1.003089e-36, -1.28498e-20, 1.027984e-20, -1.027984e-20, 
    -1.027984e-20, 1.027984e-20, -2.569961e-21, 5.139921e-21, -2.569961e-21, 
    1.003089e-36, 2.569961e-21, -5.139921e-21, -1.027984e-20, -7.709882e-21, 
    -7.709882e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, 0, 
    -1.003089e-36, 2.569961e-21, -1.541976e-20, 7.709882e-21, 1.541976e-20, 
    2.569961e-21, -2.569961e-21, -2.569961e-21, -1.003089e-36, 1.28498e-20, 
    5.139921e-21, -1.541976e-20, 2.569961e-21, 1.541976e-20, 5.139921e-21, 
    1.003089e-36, -1.003089e-36, 0, 1.027984e-20, 1.541976e-20, 
    -5.139921e-21, 5.139921e-21, 1.003089e-36, 7.709882e-21, -2.569961e-21, 
    2.569961e-21, -1.027984e-20, -1.28498e-20, -1.027984e-20, -5.139921e-21, 
    1.003089e-36, -7.709882e-21, 7.709882e-21, -1.28498e-20, -7.709882e-21, 
    5.139921e-21, 1.541976e-20, 5.139921e-21, -1.798972e-20, 2.569961e-21, 0, 
    2.569961e-21, -1.027984e-20, -7.709882e-21, -1.027984e-20, 2.569961e-21, 
    7.709882e-21, 0, 0, 2.569961e-21, -2.569961e-21, 0, -5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 1.027984e-20, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 0, 1.541976e-20, 2.569961e-21, 
    -5.139921e-21, 5.139921e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, 
    5.139921e-21, -7.709882e-21, 2.569961e-21, -1.541976e-20, -7.709882e-21, 
    -2.569961e-21, -7.709882e-21, 2.569961e-21, -2.569961e-21, 1.027984e-20, 
    1.798972e-20, -7.709882e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, 
    1.027984e-20, -7.709882e-21, 1.28498e-20, 0, 2.569961e-21, 7.709882e-21, 
    -7.709882e-21, 5.139921e-21, -1.027984e-20, 2.569961e-21, 7.709882e-21, 
    5.139921e-21, 1.027984e-20, 1.541976e-20, -2.569961e-21, -1.027984e-20, 
    -1.027984e-20, -7.709882e-21, 5.139921e-21, 5.139921e-21, -1.027984e-20, 
    2.569961e-21, -1.027984e-20, 1.027984e-20, 5.139921e-21, 2.569961e-21, 
    5.139921e-21, -1.027984e-20, 2.569961e-21, 0, 1.28498e-20, 2.569961e-21, 
    -1.027984e-20, -1.541976e-20, 2.569961e-21, -5.139921e-21, 1.027984e-20, 
    5.139921e-21, 7.709882e-21, -2.569961e-21, 0, -1.541976e-20, 
    5.139921e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, -2.569961e-21, 
    -1.003089e-36, -5.139921e-21, 1.027984e-20, -5.139921e-21, 2.569961e-21, 
    1.541976e-20, 0, 2.569961e-21, 7.709882e-21, -2.569961e-21, 
    -1.027984e-20, -1.003089e-36, -2.569961e-21, -5.139921e-21, 0, 
    -1.027984e-20, -1.541976e-20, -2.569961e-21, 5.139921e-21, -2.569961e-21, 
    5.139921e-21, 7.709882e-21, 5.139921e-21, 5.139921e-21, -2.569961e-21, 
    -5.139921e-21, 5.139921e-21, -1.798972e-20, 7.709882e-21, -2.569961e-21, 
    5.139921e-21, -7.709882e-21, -1.003089e-36, 2.569961e-21, 1.28498e-20, 
    -2.569961e-21, 5.139921e-21, -5.139921e-21, -1.28498e-20, 5.139921e-21, 
    2.569961e-21, 5.139921e-21, -2.569961e-21, -1.541976e-20, -5.139921e-21, 
    -1.28498e-20,
  1.027984e-20, 7.709882e-21, 1.027984e-20, 0, -1.027984e-20, 0, 
    -1.027984e-20, -7.709882e-21, -5.139921e-21, -7.709882e-21, 
    -7.709882e-21, 1.003089e-36, 5.139921e-21, 1.027984e-20, -5.139921e-21, 
    -7.709882e-21, 5.139921e-21, -1.027984e-20, 1.027984e-20, 1.798972e-20, 
    7.709882e-21, -1.541976e-20, -1.027984e-20, 1.027984e-20, 1.027984e-20, 
    1.027984e-20, -7.709882e-21, 1.28498e-20, 5.139921e-21, -2.569961e-21, 
    -1.003089e-36, -2.569961e-21, 1.027984e-20, -2.569961e-21, -2.569961e-21, 
    1.541976e-20, -7.709882e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    1.027984e-20, 2.569961e-21, 5.139921e-21, 1.28498e-20, 5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 0, 2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, -5.139921e-21, 1.003089e-36, 
    -7.709882e-21, -1.027984e-20, -1.027984e-20, 1.003089e-36, 7.709882e-21, 
    -7.709882e-21, 7.709882e-21, -1.28498e-20, -2.569961e-21, 1.798972e-20, 
    -7.709882e-21, 5.139921e-21, -2.055969e-20, -2.569961e-21, -5.139921e-21, 
    0, 2.569961e-21, 0, -1.027984e-20, -5.139921e-21, 1.027984e-20, 
    7.709882e-21, -2.569961e-21, 1.027984e-20, 2.569961e-21, 1.003089e-36, 
    1.28498e-20, 2.569961e-21, 1.798972e-20, -2.569961e-21, -5.139921e-21, 
    -2.312965e-20, -2.569961e-21, -7.709882e-21, -5.139921e-21, 
    -7.709882e-21, 1.003089e-36, 1.541976e-20, -1.541976e-20, -5.139921e-21, 
    -1.28498e-20, -1.027984e-20, 2.569961e-21, 1.541976e-20, -2.569961e-21, 
    -5.139921e-21, 2.055969e-20, -7.709882e-21, 7.709882e-21, -2.569961e-21, 
    1.541976e-20, -7.709882e-21, -1.027984e-20, 7.709882e-21, 7.709882e-21, 
    -1.027984e-20, 1.798972e-20, 7.709882e-21, 1.798972e-20, 7.709882e-21, 0, 
    -1.027984e-20, -1.003089e-36, -2.569961e-21, -7.709882e-21, 5.139921e-21, 
    -2.569961e-21, -7.709882e-21, -5.139921e-21, 2.569961e-20, 7.709882e-21, 
    -5.139921e-21, 5.139921e-21, -7.709882e-21, -1.027984e-20, -5.139921e-21, 
    -7.709882e-21, -1.003089e-36, 7.709882e-21, 7.709882e-21, 1.027984e-20, 
    1.027984e-20, -2.569961e-21, 0, 7.709882e-21, 5.139921e-21, 2.569961e-21, 
    -1.003089e-36, -1.027984e-20, 7.709882e-21, -2.569961e-21, -2.569961e-21, 
    -7.709882e-21, 2.569961e-21, 2.569961e-21, 0, 2.569961e-21, 1.003089e-36, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, -2.569961e-21, -2.055969e-20, 
    -5.139921e-21, 1.541976e-20, 2.569961e-21, -2.569961e-21, 1.003089e-36, 
    7.709882e-21, 7.709882e-21, -2.569961e-21, 2.569961e-21, 0, 7.709882e-21, 
    -7.709882e-21, 5.139921e-21, -1.28498e-20, 5.139921e-21, -1.541976e-20, 
    0, 1.28498e-20, 2.569961e-21, -7.709882e-21, 5.139921e-21, 1.003089e-36, 
    1.027984e-20, 0, -5.139921e-21, -5.139921e-21, 1.798972e-20, 
    -1.027984e-20, -7.709882e-21, 1.027984e-20, 2.569961e-21, 7.709882e-21, 
    -1.027984e-20, 2.569961e-21, 2.569961e-21, -7.709882e-21, 1.003089e-36, 
    0, 2.569961e-21, -1.027984e-20, -5.139921e-21, -2.569961e-21, 
    -5.139921e-21, 0, 1.027984e-20, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, 0, 2.569961e-21, -2.055969e-20, -1.28498e-20, 
    -2.569961e-21, 0, -7.709882e-21, 5.139921e-21, -1.28498e-20, 
    -2.569961e-21, 5.139921e-21, 7.709882e-21, 1.798972e-20, 1.798972e-20, 
    -5.139921e-21, -2.569961e-21, -1.027984e-20, -7.709882e-21, 1.027984e-20, 
    2.569961e-21, 1.541976e-20, -2.569961e-21, 2.569961e-21, -1.027984e-20, 
    -2.569961e-21, -7.709882e-21, -7.709882e-21, 0, 2.569961e-21, 
    5.139921e-21, 1.003089e-36, 5.139921e-21, -7.709882e-21, -1.003089e-36, 
    1.027984e-20, -1.28498e-20, 5.139921e-21, -1.027984e-20, 7.709882e-21, 
    2.569961e-21, 2.569961e-21, 2.569961e-21, 5.139921e-21, -5.139921e-21, 
    7.709882e-21, 1.28498e-20, 2.569961e-21, -5.139921e-21, -1.003089e-36, 
    -7.709882e-21, 1.027984e-20, -1.027984e-20, 5.139921e-21, 5.139921e-21, 
    2.055969e-20, -5.139921e-21, -7.709882e-21, -1.28498e-20, -2.569961e-21, 
    -7.709882e-21, 1.027984e-20, -1.28498e-20, -2.055969e-20, 2.055969e-20, 
    -2.055969e-20, 5.139921e-21, -7.709882e-21, 0, -1.541976e-20, 
    -1.003089e-36, -2.055969e-20, 0, -5.139921e-21, -7.709882e-21, 
    -5.139921e-21, 5.139921e-21, -1.003089e-36, 7.709882e-21, -5.139921e-21, 
    -2.569961e-21, 5.139921e-21, -1.798972e-20, 2.569961e-21, -2.569961e-21, 
    5.139921e-21, -2.569961e-21, -7.709882e-21, 2.569961e-21, -7.709882e-21, 
    1.28498e-20, 2.569961e-21, 1.28498e-20, -1.027984e-20, -5.139921e-21, 
    5.139921e-21, -1.027984e-20, 0, 1.28498e-20, -5.139921e-21, 2.569961e-21, 
    5.139921e-21, -2.569961e-21, -1.798972e-20, 1.027984e-20, 1.798972e-20, 
    -7.709882e-21, 2.569961e-21, -2.055969e-20, 1.28498e-20, -2.569961e-21, 
    -1.28498e-20, 7.709882e-21, -1.541976e-20, -1.28498e-20, -5.139921e-21, 
    -2.569961e-21, 2.569961e-21, -7.709882e-21, -7.709882e-21, -7.709882e-21, 
    -2.569961e-21, -1.798972e-20, 1.027984e-20, 7.709882e-21, 5.139921e-21, 
    -5.139921e-21, -7.709882e-21, 5.139921e-21, 5.139921e-21, -1.027984e-20, 
    -5.139921e-21, -5.139921e-21,
  5.139921e-21, 0, 1.027984e-20, 1.28498e-20, -7.709882e-21, -5.139921e-21, 
    -1.798972e-20, -2.312965e-20, 5.139921e-21, 2.055969e-20, -1.003089e-36, 
    -1.027984e-20, -7.709882e-21, -1.027984e-20, 1.027984e-20, -1.027984e-20, 
    -7.709882e-21, 5.139921e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, 
    1.003089e-36, 2.569961e-21, -7.709882e-21, 2.312965e-20, -3.083953e-20, 
    5.139921e-21, -2.569961e-21, -7.709882e-21, 2.055969e-20, -1.541976e-20, 
    -2.569961e-21, -2.569961e-21, -1.541976e-20, -2.569961e-21, 7.709882e-21, 
    2.569961e-21, 1.28498e-20, 2.569961e-21, 5.139921e-21, -1.28498e-20, 
    7.709882e-21, -1.027984e-20, -2.312965e-20, -1.003089e-36, -2.569961e-21, 
    -1.541976e-20, 5.139921e-21, 2.569961e-21, 7.709882e-21, -2.569961e-21, 
    2.055969e-20, 0, 1.027984e-20, -5.139921e-21, -2.826957e-20, 
    -1.541976e-20, 7.709882e-21, -1.28498e-20, 1.28498e-20, 1.28498e-20, 
    1.003089e-36, 7.709882e-21, 2.569961e-21, -1.28498e-20, 5.139921e-21, 
    5.139921e-21, -2.312965e-20, -5.139921e-21, -1.798972e-20, -7.709882e-21, 
    1.027984e-20, 2.569961e-21, -2.569961e-21, 1.027984e-20, 1.541976e-20, 
    -2.569961e-21, 1.027984e-20, -7.709882e-21, -2.569961e-21, 1.027984e-20, 
    7.709882e-21, 5.139921e-21, 2.569961e-21, 7.709882e-21, -2.569961e-21, 
    7.709882e-21, 1.28498e-20, 1.541976e-20, 2.055969e-20, -2.569961e-21, 
    -2.055969e-20, 1.798972e-20, 1.28498e-20, -7.709882e-21, -5.139921e-21, 
    -1.027984e-20, 1.003089e-36, 2.569961e-21, 1.003089e-36, -1.541976e-20, 
    -1.28498e-20, -1.28498e-20, 5.139921e-21, -7.709882e-21, 1.027984e-20, 
    -1.027984e-20, 1.027984e-20, -1.28498e-20, -2.569961e-21, 1.28498e-20, 
    -2.055969e-20, 1.027984e-20, 2.569961e-21, 1.28498e-20, -7.709882e-21, 
    7.709882e-21, 1.003089e-36, 2.569961e-21, -2.055969e-20, -2.055969e-20, 
    -1.28498e-20, -1.798972e-20, 1.28498e-20, 2.312965e-20, 5.139921e-21, 
    1.798972e-20, 1.003089e-36, 1.027984e-20, 1.541976e-20, -1.027984e-20, 
    -2.569961e-21, -5.139921e-21, 2.055969e-20, 1.28498e-20, -1.28498e-20, 
    1.027984e-20, 1.027984e-20, -1.027984e-20, -7.709882e-21, -2.569961e-21, 
    1.027984e-20, -7.709882e-21, 2.312965e-20, -1.28498e-20, -2.312965e-20, 
    -1.027984e-20, -1.027984e-20, -5.139921e-21, 2.569961e-21, -1.541976e-20, 
    2.569961e-21, 1.027984e-20, -5.139921e-21, 2.569961e-21, 1.541976e-20, 
    -2.569961e-21, 2.569961e-21, -7.709882e-21, -2.569961e-21, -7.709882e-21, 
    -2.569961e-21, -1.003089e-36, -3.340949e-20, -1.28498e-20, -1.28498e-20, 
    -7.709882e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, -7.709882e-21, 
    1.798972e-20, 5.139921e-21, 3.597945e-20, -1.798972e-20, -5.139921e-21, 
    7.709882e-21, 1.28498e-20, 7.709882e-21, -1.798972e-20, 7.709882e-21, 
    5.139921e-21, -2.569961e-21, 5.139921e-21, -1.541976e-20, -2.569961e-21, 
    7.709882e-21, -1.541976e-20, -7.709882e-21, -1.28498e-20, -1.027984e-20, 
    2.569961e-21, 1.003089e-36, 2.569961e-21, 1.027984e-20, 7.709882e-21, 
    7.709882e-21, 7.709882e-21, 0, -5.139921e-21, -1.28498e-20, 2.569961e-21, 
    1.541976e-20, -2.312965e-20, -2.569961e-21, 5.139921e-21, -1.003089e-36, 
    -2.569961e-21, -1.28498e-20, 1.798972e-20, -7.709882e-21, -1.541976e-20, 
    1.027984e-20, 2.055969e-20, -2.569961e-21, -2.569961e-21, 2.569961e-21, 
    -1.28498e-20, -2.826957e-20, -1.003089e-36, -1.027984e-20, 1.541976e-20, 
    7.709882e-21, 2.569961e-21, 2.569961e-21, -7.709882e-21, 3.083953e-20, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, 5.139921e-21, 1.541976e-20, 
    5.139921e-21, -1.28498e-20, -5.139921e-21, -7.709882e-21, -5.139921e-21, 
    -7.709882e-21, 1.28498e-20, 7.709882e-21, -1.28498e-20, 1.027984e-20, 
    2.055969e-20, 1.28498e-20, 1.027984e-20, 1.541976e-20, -2.826957e-20, 
    -5.139921e-21, 1.28498e-20, 2.569961e-21, 7.709882e-21, 1.027984e-20, 
    -1.027984e-20, -5.139921e-21, 0, 7.709882e-21, 7.709882e-21, 
    1.541976e-20, -7.709882e-21, -7.709882e-21, -7.709882e-21, -1.28498e-20, 
    1.798972e-20, -7.709882e-21, -1.027984e-20, 1.027984e-20, -2.312965e-20, 
    2.569961e-21, 2.569961e-21, -2.569961e-21, -1.027984e-20, -2.569961e-21, 
    -2.569961e-21, -2.569961e-21, 5.139921e-21, 0, 2.569961e-21, 0, 
    2.055969e-20, 2.569961e-21, 7.709882e-21, -2.569961e-21, -7.709882e-21, 
    2.569961e-21, 5.139921e-21, 7.709882e-21, -2.569961e-21, 2.569961e-21, 
    -1.541976e-20, 2.569961e-21, 0, -5.139921e-21, -1.28498e-20, 
    -1.541976e-20, 3.340949e-20, -1.027984e-20, 1.28498e-20, -5.139921e-21, 
    -5.139921e-21, 2.569961e-21, -7.709882e-21, 1.798972e-20, -1.003089e-36, 
    -5.139921e-21, -1.027984e-20, -7.709882e-21, 7.709882e-21, -1.027984e-20, 
    1.027984e-20, 5.139921e-21, -1.027984e-20, -5.139921e-21, -2.569961e-20, 
    -1.003089e-36, 1.541976e-20, -5.139921e-21, -7.709882e-21, -5.139921e-21, 
    7.709882e-21, -1.003089e-36, 5.139921e-21, 7.709882e-21, 1.28498e-20, 
    -7.709882e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, 2.006177e-36, 
    -2.569961e-21, -1.027984e-20, -1.027984e-20, -5.139921e-21, 2.569961e-21, 
    -1.003089e-36, -5.139921e-21, 0, -2.569961e-21, -1.027984e-20,
  6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N_TO_SOIL1N =
  5.288484e-12, 5.311751e-12, 5.307228e-12, 5.325994e-12, 5.315583e-12, 
    5.327872e-12, 5.293201e-12, 5.312675e-12, 5.300243e-12, 5.290578e-12, 
    5.362413e-12, 5.326831e-12, 5.39937e-12, 5.376678e-12, 5.43368e-12, 
    5.395839e-12, 5.44131e-12, 5.432588e-12, 5.458838e-12, 5.451318e-12, 
    5.484896e-12, 5.462309e-12, 5.5023e-12, 5.479501e-12, 5.483068e-12, 
    5.461564e-12, 5.333991e-12, 5.357983e-12, 5.332569e-12, 5.335991e-12, 
    5.334456e-12, 5.315799e-12, 5.306397e-12, 5.286706e-12, 5.29028e-12, 
    5.304743e-12, 5.337529e-12, 5.326399e-12, 5.354448e-12, 5.353815e-12, 
    5.385041e-12, 5.370961e-12, 5.423444e-12, 5.408528e-12, 5.451632e-12, 
    5.440792e-12, 5.451123e-12, 5.44799e-12, 5.451163e-12, 5.435265e-12, 
    5.442077e-12, 5.428087e-12, 5.373598e-12, 5.389612e-12, 5.341851e-12, 
    5.313132e-12, 5.294055e-12, 5.280519e-12, 5.282432e-12, 5.286081e-12, 
    5.304828e-12, 5.322453e-12, 5.335885e-12, 5.34487e-12, 5.353724e-12, 
    5.380522e-12, 5.394704e-12, 5.426461e-12, 5.420729e-12, 5.430439e-12, 
    5.439713e-12, 5.455286e-12, 5.452722e-12, 5.459583e-12, 5.430182e-12, 
    5.449722e-12, 5.417465e-12, 5.426287e-12, 5.356133e-12, 5.329402e-12, 
    5.318042e-12, 5.308097e-12, 5.283904e-12, 5.300612e-12, 5.294025e-12, 
    5.309694e-12, 5.31965e-12, 5.314726e-12, 5.345116e-12, 5.333301e-12, 
    5.395545e-12, 5.368735e-12, 5.438631e-12, 5.421906e-12, 5.44264e-12, 
    5.43206e-12, 5.450189e-12, 5.433873e-12, 5.462136e-12, 5.468291e-12, 
    5.464085e-12, 5.48024e-12, 5.432968e-12, 5.451123e-12, 5.314588e-12, 
    5.315391e-12, 5.319132e-12, 5.302686e-12, 5.30168e-12, 5.286608e-12, 
    5.300019e-12, 5.30573e-12, 5.320227e-12, 5.328802e-12, 5.336954e-12, 
    5.354877e-12, 5.374893e-12, 5.402882e-12, 5.42299e-12, 5.436469e-12, 
    5.428203e-12, 5.4355e-12, 5.427343e-12, 5.42352e-12, 5.465985e-12, 
    5.442141e-12, 5.477917e-12, 5.475937e-12, 5.459746e-12, 5.47616e-12, 
    5.315955e-12, 5.311333e-12, 5.295288e-12, 5.307845e-12, 5.284966e-12, 
    5.297773e-12, 5.305137e-12, 5.333549e-12, 5.33979e-12, 5.345579e-12, 
    5.357011e-12, 5.371682e-12, 5.397419e-12, 5.419811e-12, 5.440253e-12, 
    5.438755e-12, 5.439282e-12, 5.443849e-12, 5.432537e-12, 5.445706e-12, 
    5.447916e-12, 5.442138e-12, 5.475672e-12, 5.466092e-12, 5.475895e-12, 
    5.469657e-12, 5.312835e-12, 5.320612e-12, 5.31641e-12, 5.324312e-12, 
    5.318745e-12, 5.343498e-12, 5.35092e-12, 5.385645e-12, 5.371393e-12, 
    5.394075e-12, 5.373697e-12, 5.377308e-12, 5.394816e-12, 5.374798e-12, 
    5.418577e-12, 5.388897e-12, 5.444027e-12, 5.414389e-12, 5.445884e-12, 
    5.440164e-12, 5.449634e-12, 5.458115e-12, 5.468784e-12, 5.488471e-12, 
    5.483912e-12, 5.500375e-12, 5.332205e-12, 5.342291e-12, 5.341403e-12, 
    5.351958e-12, 5.359764e-12, 5.376683e-12, 5.403819e-12, 5.393615e-12, 
    5.412348e-12, 5.416109e-12, 5.387648e-12, 5.405123e-12, 5.349041e-12, 
    5.358103e-12, 5.352707e-12, 5.333001e-12, 5.395967e-12, 5.363653e-12, 
    5.423322e-12, 5.405817e-12, 5.456906e-12, 5.431499e-12, 5.481403e-12, 
    5.502737e-12, 5.522814e-12, 5.546279e-12, 5.347796e-12, 5.340942e-12, 
    5.353213e-12, 5.370191e-12, 5.385943e-12, 5.406885e-12, 5.409027e-12, 
    5.41295e-12, 5.423112e-12, 5.431657e-12, 5.414192e-12, 5.433798e-12, 
    5.360205e-12, 5.398772e-12, 5.338351e-12, 5.356546e-12, 5.36919e-12, 
    5.363643e-12, 5.392449e-12, 5.399238e-12, 5.426827e-12, 5.412564e-12, 
    5.497472e-12, 5.459907e-12, 5.564143e-12, 5.535014e-12, 5.338547e-12, 
    5.347772e-12, 5.379875e-12, 5.3646e-12, 5.408283e-12, 5.419035e-12, 
    5.427775e-12, 5.438949e-12, 5.440155e-12, 5.446775e-12, 5.435927e-12, 
    5.446347e-12, 5.406929e-12, 5.424544e-12, 5.376205e-12, 5.387971e-12, 
    5.382558e-12, 5.376621e-12, 5.394944e-12, 5.414467e-12, 5.414883e-12, 
    5.421143e-12, 5.438784e-12, 5.40846e-12, 5.502322e-12, 5.444356e-12, 
    5.35783e-12, 5.375598e-12, 5.378135e-12, 5.371252e-12, 5.417957e-12, 
    5.401034e-12, 5.446614e-12, 5.434295e-12, 5.454479e-12, 5.44445e-12, 
    5.442974e-12, 5.430092e-12, 5.422072e-12, 5.401811e-12, 5.385324e-12, 
    5.37225e-12, 5.37529e-12, 5.389651e-12, 5.415661e-12, 5.440265e-12, 
    5.434875e-12, 5.452945e-12, 5.405115e-12, 5.425172e-12, 5.41742e-12, 
    5.437632e-12, 5.393344e-12, 5.43106e-12, 5.383703e-12, 5.387856e-12, 
    5.400699e-12, 5.426532e-12, 5.432247e-12, 5.43835e-12, 5.434584e-12, 
    5.416321e-12, 5.413328e-12, 5.400386e-12, 5.396813e-12, 5.386951e-12, 
    5.378787e-12, 5.386247e-12, 5.394081e-12, 5.416328e-12, 5.436377e-12, 
    5.458235e-12, 5.463584e-12, 5.489126e-12, 5.468335e-12, 5.502645e-12, 
    5.473477e-12, 5.523967e-12, 5.433244e-12, 5.472618e-12, 5.401283e-12, 
    5.408968e-12, 5.422868e-12, 5.454749e-12, 5.437537e-12, 5.457666e-12, 
    5.413211e-12, 5.390148e-12, 5.384179e-12, 5.373045e-12, 5.384434e-12, 
    5.383507e-12, 5.394405e-12, 5.390903e-12, 5.417067e-12, 5.403013e-12, 
    5.442937e-12, 5.457506e-12, 5.49865e-12, 5.523873e-12, 5.549547e-12, 
    5.560882e-12, 5.564332e-12, 5.565774e-12 ;

 SOIL3N_vr =
  1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.81819, 1.81819, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.81819, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818188, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3_HR =
  3.199533e-11, 3.213609e-11, 3.210873e-11, 3.222226e-11, 3.215928e-11, 
    3.223363e-11, 3.202387e-11, 3.214168e-11, 3.206647e-11, 3.2008e-11, 
    3.24426e-11, 3.222733e-11, 3.266619e-11, 3.25289e-11, 3.287377e-11, 
    3.264482e-11, 3.291993e-11, 3.286716e-11, 3.302597e-11, 3.298047e-11, 
    3.318362e-11, 3.304697e-11, 3.328891e-11, 3.315098e-11, 3.317256e-11, 
    3.304246e-11, 3.227064e-11, 3.24158e-11, 3.226205e-11, 3.228275e-11, 
    3.227345e-11, 3.216058e-11, 3.210371e-11, 3.198457e-11, 3.20062e-11, 
    3.20937e-11, 3.229205e-11, 3.222472e-11, 3.239441e-11, 3.239058e-11, 
    3.257949e-11, 3.249432e-11, 3.281184e-11, 3.272159e-11, 3.298237e-11, 
    3.291679e-11, 3.297929e-11, 3.296034e-11, 3.297954e-11, 3.288336e-11, 
    3.292457e-11, 3.283993e-11, 3.251027e-11, 3.260716e-11, 3.23182e-11, 
    3.214445e-11, 3.202904e-11, 3.194714e-11, 3.195871e-11, 3.198079e-11, 
    3.209421e-11, 3.220084e-11, 3.228211e-11, 3.233647e-11, 3.239003e-11, 
    3.255216e-11, 3.263796e-11, 3.283009e-11, 3.279541e-11, 3.285415e-11, 
    3.291026e-11, 3.300448e-11, 3.298897e-11, 3.303048e-11, 3.28526e-11, 
    3.297082e-11, 3.277566e-11, 3.282904e-11, 3.24046e-11, 3.224288e-11, 
    3.217416e-11, 3.211399e-11, 3.196762e-11, 3.20687e-11, 3.202885e-11, 
    3.212365e-11, 3.218388e-11, 3.215409e-11, 3.233795e-11, 3.226647e-11, 
    3.264305e-11, 3.248084e-11, 3.290372e-11, 3.280253e-11, 3.292797e-11, 
    3.286396e-11, 3.297364e-11, 3.287493e-11, 3.304593e-11, 3.308316e-11, 
    3.305772e-11, 3.315545e-11, 3.286946e-11, 3.297929e-11, 3.215326e-11, 
    3.215811e-11, 3.218075e-11, 3.208125e-11, 3.207516e-11, 3.198397e-11, 
    3.206511e-11, 3.209967e-11, 3.218737e-11, 3.223925e-11, 3.228857e-11, 
    3.239701e-11, 3.25181e-11, 3.268744e-11, 3.280909e-11, 3.289063e-11, 
    3.284063e-11, 3.288478e-11, 3.283543e-11, 3.281229e-11, 3.306921e-11, 
    3.292495e-11, 3.31414e-11, 3.312942e-11, 3.303147e-11, 3.313077e-11, 
    3.216153e-11, 3.213357e-11, 3.203649e-11, 3.211246e-11, 3.197404e-11, 
    3.205152e-11, 3.209608e-11, 3.226797e-11, 3.230573e-11, 3.234075e-11, 
    3.240992e-11, 3.249868e-11, 3.265438e-11, 3.278986e-11, 3.291353e-11, 
    3.290447e-11, 3.290766e-11, 3.293529e-11, 3.286685e-11, 3.294652e-11, 
    3.29599e-11, 3.292493e-11, 3.312782e-11, 3.306985e-11, 3.312917e-11, 
    3.309143e-11, 3.214265e-11, 3.21897e-11, 3.216428e-11, 3.221208e-11, 
    3.217841e-11, 3.232816e-11, 3.237306e-11, 3.258315e-11, 3.249693e-11, 
    3.263415e-11, 3.251087e-11, 3.253271e-11, 3.263863e-11, 3.251753e-11, 
    3.278239e-11, 3.260283e-11, 3.293636e-11, 3.275705e-11, 3.29476e-11, 
    3.2913e-11, 3.297028e-11, 3.30216e-11, 3.308614e-11, 3.320525e-11, 
    3.317767e-11, 3.327727e-11, 3.225984e-11, 3.232086e-11, 3.231549e-11, 
    3.237935e-11, 3.242657e-11, 3.252893e-11, 3.269311e-11, 3.263137e-11, 
    3.274471e-11, 3.276746e-11, 3.259527e-11, 3.270099e-11, 3.23617e-11, 
    3.241652e-11, 3.238388e-11, 3.226465e-11, 3.26456e-11, 3.24501e-11, 
    3.28111e-11, 3.270519e-11, 3.301428e-11, 3.286057e-11, 3.316248e-11, 
    3.329156e-11, 3.341302e-11, 3.355499e-11, 3.235416e-11, 3.23127e-11, 
    3.238694e-11, 3.248966e-11, 3.258496e-11, 3.271165e-11, 3.272461e-11, 
    3.274835e-11, 3.280983e-11, 3.286152e-11, 3.275586e-11, 3.287448e-11, 
    3.242924e-11, 3.266257e-11, 3.229703e-11, 3.24071e-11, 3.24836e-11, 
    3.245004e-11, 3.262431e-11, 3.266539e-11, 3.28323e-11, 3.274601e-11, 
    3.32597e-11, 3.303243e-11, 3.366307e-11, 3.348683e-11, 3.229821e-11, 
    3.235402e-11, 3.254825e-11, 3.245583e-11, 3.272011e-11, 3.278516e-11, 
    3.283804e-11, 3.290564e-11, 3.291294e-11, 3.295299e-11, 3.288736e-11, 
    3.29504e-11, 3.271192e-11, 3.281849e-11, 3.252604e-11, 3.259722e-11, 
    3.256448e-11, 3.252856e-11, 3.263942e-11, 3.275752e-11, 3.276004e-11, 
    3.279791e-11, 3.290464e-11, 3.272118e-11, 3.328905e-11, 3.293835e-11, 
    3.241487e-11, 3.252237e-11, 3.253772e-11, 3.249608e-11, 3.277864e-11, 
    3.267626e-11, 3.295202e-11, 3.287749e-11, 3.29996e-11, 3.293892e-11, 
    3.292999e-11, 3.285206e-11, 3.280354e-11, 3.268096e-11, 3.258121e-11, 
    3.250212e-11, 3.252051e-11, 3.260739e-11, 3.276475e-11, 3.29136e-11, 
    3.288099e-11, 3.299032e-11, 3.270095e-11, 3.282229e-11, 3.277539e-11, 
    3.289767e-11, 3.262973e-11, 3.285791e-11, 3.257141e-11, 3.259653e-11, 
    3.267422e-11, 3.283052e-11, 3.286509e-11, 3.290201e-11, 3.287923e-11, 
    3.276874e-11, 3.275064e-11, 3.267234e-11, 3.265072e-11, 3.259105e-11, 
    3.254166e-11, 3.258679e-11, 3.263419e-11, 3.276878e-11, 3.289008e-11, 
    3.302232e-11, 3.305469e-11, 3.320921e-11, 3.308343e-11, 3.3291e-11, 
    3.311454e-11, 3.342e-11, 3.287113e-11, 3.310933e-11, 3.267776e-11, 
    3.272425e-11, 3.280835e-11, 3.300123e-11, 3.28971e-11, 3.301888e-11, 
    3.274993e-11, 3.261039e-11, 3.257428e-11, 3.250692e-11, 3.257582e-11, 
    3.257022e-11, 3.263615e-11, 3.261496e-11, 3.277325e-11, 3.268823e-11, 
    3.292977e-11, 3.301791e-11, 3.326683e-11, 3.341943e-11, 3.357476e-11, 
    3.364333e-11, 3.366421e-11, 3.367293e-11 ;

 SOILC =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34457, 17.34459, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.3446, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34456, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34452, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.3445, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.34449, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34457, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34453, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34456, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34455, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 SOILC_HR =
  6.357484e-08, 6.385439e-08, 6.380004e-08, 6.402553e-08, 6.390044e-08, 
    6.404809e-08, 6.363151e-08, 6.386549e-08, 6.371612e-08, 6.360001e-08, 
    6.446311e-08, 6.403558e-08, 6.490716e-08, 6.463451e-08, 6.53194e-08, 
    6.486474e-08, 6.541108e-08, 6.530627e-08, 6.562168e-08, 6.553132e-08, 
    6.593476e-08, 6.566339e-08, 6.614388e-08, 6.586995e-08, 6.59128e-08, 
    6.565443e-08, 6.412161e-08, 6.440989e-08, 6.410454e-08, 6.414565e-08, 
    6.41272e-08, 6.390303e-08, 6.379007e-08, 6.355347e-08, 6.359642e-08, 
    6.377019e-08, 6.416413e-08, 6.40304e-08, 6.436741e-08, 6.43598e-08, 
    6.473498e-08, 6.456582e-08, 6.519642e-08, 6.501719e-08, 6.55351e-08, 
    6.540485e-08, 6.552898e-08, 6.549134e-08, 6.552947e-08, 6.533845e-08, 
    6.542029e-08, 6.52522e-08, 6.459751e-08, 6.478992e-08, 6.421605e-08, 
    6.387099e-08, 6.364178e-08, 6.347913e-08, 6.350213e-08, 6.354596e-08, 
    6.377121e-08, 6.398299e-08, 6.414438e-08, 6.425233e-08, 6.43587e-08, 
    6.46807e-08, 6.48511e-08, 6.523266e-08, 6.51638e-08, 6.528045e-08, 
    6.539189e-08, 6.557899e-08, 6.55482e-08, 6.563063e-08, 6.527737e-08, 
    6.551215e-08, 6.512457e-08, 6.523057e-08, 6.438765e-08, 6.406648e-08, 
    6.392999e-08, 6.38105e-08, 6.351981e-08, 6.372055e-08, 6.364142e-08, 
    6.382967e-08, 6.39493e-08, 6.389013e-08, 6.425529e-08, 6.411333e-08, 
    6.48612e-08, 6.453907e-08, 6.537889e-08, 6.517793e-08, 6.542706e-08, 
    6.529993e-08, 6.551776e-08, 6.532171e-08, 6.566131e-08, 6.573526e-08, 
    6.568472e-08, 6.587883e-08, 6.531085e-08, 6.552898e-08, 6.388848e-08, 
    6.389813e-08, 6.394308e-08, 6.374548e-08, 6.373339e-08, 6.355229e-08, 
    6.371343e-08, 6.378205e-08, 6.395624e-08, 6.405927e-08, 6.415721e-08, 
    6.437256e-08, 6.461306e-08, 6.494936e-08, 6.519095e-08, 6.53529e-08, 
    6.525359e-08, 6.534127e-08, 6.524326e-08, 6.519733e-08, 6.570755e-08, 
    6.542106e-08, 6.585091e-08, 6.582712e-08, 6.563259e-08, 6.582981e-08, 
    6.390491e-08, 6.384938e-08, 6.365659e-08, 6.380746e-08, 6.353257e-08, 
    6.368644e-08, 6.377493e-08, 6.41163e-08, 6.41913e-08, 6.426085e-08, 
    6.43982e-08, 6.457448e-08, 6.488371e-08, 6.515276e-08, 6.539837e-08, 
    6.538038e-08, 6.538671e-08, 6.544158e-08, 6.530567e-08, 6.546389e-08, 
    6.549045e-08, 6.542102e-08, 6.582394e-08, 6.570883e-08, 6.582662e-08, 
    6.575167e-08, 6.386743e-08, 6.396086e-08, 6.391037e-08, 6.400531e-08, 
    6.393843e-08, 6.423585e-08, 6.432501e-08, 6.474225e-08, 6.457101e-08, 
    6.484353e-08, 6.459869e-08, 6.464208e-08, 6.485244e-08, 6.461192e-08, 
    6.513793e-08, 6.478133e-08, 6.544371e-08, 6.508762e-08, 6.546603e-08, 
    6.539731e-08, 6.551109e-08, 6.561299e-08, 6.574118e-08, 6.597772e-08, 
    6.592295e-08, 6.612076e-08, 6.410015e-08, 6.422135e-08, 6.421067e-08, 
    6.433749e-08, 6.443128e-08, 6.463457e-08, 6.496062e-08, 6.483801e-08, 
    6.506309e-08, 6.510828e-08, 6.476632e-08, 6.497628e-08, 6.430245e-08, 
    6.441132e-08, 6.434649e-08, 6.410971e-08, 6.486627e-08, 6.447801e-08, 
    6.519495e-08, 6.498462e-08, 6.559846e-08, 6.529319e-08, 6.589279e-08, 
    6.614913e-08, 6.639036e-08, 6.667229e-08, 6.428748e-08, 6.420513e-08, 
    6.435257e-08, 6.455657e-08, 6.474583e-08, 6.499745e-08, 6.502319e-08, 
    6.507033e-08, 6.519242e-08, 6.529509e-08, 6.508524e-08, 6.532083e-08, 
    6.443658e-08, 6.489997e-08, 6.4174e-08, 6.439262e-08, 6.454454e-08, 
    6.44779e-08, 6.482399e-08, 6.490557e-08, 6.523705e-08, 6.506569e-08, 
    6.608587e-08, 6.563452e-08, 6.688694e-08, 6.653695e-08, 6.417636e-08, 
    6.428719e-08, 6.467292e-08, 6.448939e-08, 6.501424e-08, 6.514343e-08, 
    6.524845e-08, 6.538271e-08, 6.53972e-08, 6.547674e-08, 6.53464e-08, 
    6.547159e-08, 6.499798e-08, 6.520963e-08, 6.462883e-08, 6.47702e-08, 
    6.470516e-08, 6.463382e-08, 6.485399e-08, 6.508855e-08, 6.509355e-08, 
    6.516876e-08, 6.538072e-08, 6.501637e-08, 6.614414e-08, 6.544767e-08, 
    6.440805e-08, 6.462153e-08, 6.465201e-08, 6.456932e-08, 6.513049e-08, 
    6.492716e-08, 6.54748e-08, 6.532679e-08, 6.55693e-08, 6.544879e-08, 
    6.543107e-08, 6.527629e-08, 6.517993e-08, 6.493648e-08, 6.473839e-08, 
    6.458131e-08, 6.461784e-08, 6.479039e-08, 6.51029e-08, 6.539852e-08, 
    6.533376e-08, 6.555087e-08, 6.497619e-08, 6.521717e-08, 6.512403e-08, 
    6.536688e-08, 6.483475e-08, 6.528791e-08, 6.471893e-08, 6.476881e-08, 
    6.492312e-08, 6.523352e-08, 6.530218e-08, 6.537551e-08, 6.533025e-08, 
    6.511083e-08, 6.507487e-08, 6.491937e-08, 6.487644e-08, 6.475795e-08, 
    6.465985e-08, 6.474948e-08, 6.48436e-08, 6.511091e-08, 6.535181e-08, 
    6.561444e-08, 6.567871e-08, 6.598559e-08, 6.573579e-08, 6.614802e-08, 
    6.579756e-08, 6.640422e-08, 6.531416e-08, 6.578724e-08, 6.493014e-08, 
    6.502248e-08, 6.518949e-08, 6.557254e-08, 6.536574e-08, 6.560759e-08, 
    6.507346e-08, 6.479635e-08, 6.472464e-08, 6.459086e-08, 6.472769e-08, 
    6.471657e-08, 6.48475e-08, 6.480542e-08, 6.511979e-08, 6.495092e-08, 
    6.543063e-08, 6.560568e-08, 6.610003e-08, 6.640308e-08, 6.671156e-08, 
    6.684775e-08, 6.68892e-08, 6.690653e-08 ;

 SOILC_LOSS =
  6.357484e-08, 6.385439e-08, 6.380004e-08, 6.402553e-08, 6.390044e-08, 
    6.404809e-08, 6.363151e-08, 6.386549e-08, 6.371612e-08, 6.360001e-08, 
    6.446311e-08, 6.403558e-08, 6.490716e-08, 6.463451e-08, 6.53194e-08, 
    6.486474e-08, 6.541108e-08, 6.530627e-08, 6.562168e-08, 6.553132e-08, 
    6.593476e-08, 6.566339e-08, 6.614388e-08, 6.586995e-08, 6.59128e-08, 
    6.565443e-08, 6.412161e-08, 6.440989e-08, 6.410454e-08, 6.414565e-08, 
    6.41272e-08, 6.390303e-08, 6.379007e-08, 6.355347e-08, 6.359642e-08, 
    6.377019e-08, 6.416413e-08, 6.40304e-08, 6.436741e-08, 6.43598e-08, 
    6.473498e-08, 6.456582e-08, 6.519642e-08, 6.501719e-08, 6.55351e-08, 
    6.540485e-08, 6.552898e-08, 6.549134e-08, 6.552947e-08, 6.533845e-08, 
    6.542029e-08, 6.52522e-08, 6.459751e-08, 6.478992e-08, 6.421605e-08, 
    6.387099e-08, 6.364178e-08, 6.347913e-08, 6.350213e-08, 6.354596e-08, 
    6.377121e-08, 6.398299e-08, 6.414438e-08, 6.425233e-08, 6.43587e-08, 
    6.46807e-08, 6.48511e-08, 6.523266e-08, 6.51638e-08, 6.528045e-08, 
    6.539189e-08, 6.557899e-08, 6.55482e-08, 6.563063e-08, 6.527737e-08, 
    6.551215e-08, 6.512457e-08, 6.523057e-08, 6.438765e-08, 6.406648e-08, 
    6.392999e-08, 6.38105e-08, 6.351981e-08, 6.372055e-08, 6.364142e-08, 
    6.382967e-08, 6.39493e-08, 6.389013e-08, 6.425529e-08, 6.411333e-08, 
    6.48612e-08, 6.453907e-08, 6.537889e-08, 6.517793e-08, 6.542706e-08, 
    6.529993e-08, 6.551776e-08, 6.532171e-08, 6.566131e-08, 6.573526e-08, 
    6.568472e-08, 6.587883e-08, 6.531085e-08, 6.552898e-08, 6.388848e-08, 
    6.389813e-08, 6.394308e-08, 6.374548e-08, 6.373339e-08, 6.355229e-08, 
    6.371343e-08, 6.378205e-08, 6.395624e-08, 6.405927e-08, 6.415721e-08, 
    6.437256e-08, 6.461306e-08, 6.494936e-08, 6.519095e-08, 6.53529e-08, 
    6.525359e-08, 6.534127e-08, 6.524326e-08, 6.519733e-08, 6.570755e-08, 
    6.542106e-08, 6.585091e-08, 6.582712e-08, 6.563259e-08, 6.582981e-08, 
    6.390491e-08, 6.384938e-08, 6.365659e-08, 6.380746e-08, 6.353257e-08, 
    6.368644e-08, 6.377493e-08, 6.41163e-08, 6.41913e-08, 6.426085e-08, 
    6.43982e-08, 6.457448e-08, 6.488371e-08, 6.515276e-08, 6.539837e-08, 
    6.538038e-08, 6.538671e-08, 6.544158e-08, 6.530567e-08, 6.546389e-08, 
    6.549045e-08, 6.542102e-08, 6.582394e-08, 6.570883e-08, 6.582662e-08, 
    6.575167e-08, 6.386743e-08, 6.396086e-08, 6.391037e-08, 6.400531e-08, 
    6.393843e-08, 6.423585e-08, 6.432501e-08, 6.474225e-08, 6.457101e-08, 
    6.484353e-08, 6.459869e-08, 6.464208e-08, 6.485244e-08, 6.461192e-08, 
    6.513793e-08, 6.478133e-08, 6.544371e-08, 6.508762e-08, 6.546603e-08, 
    6.539731e-08, 6.551109e-08, 6.561299e-08, 6.574118e-08, 6.597772e-08, 
    6.592295e-08, 6.612076e-08, 6.410015e-08, 6.422135e-08, 6.421067e-08, 
    6.433749e-08, 6.443128e-08, 6.463457e-08, 6.496062e-08, 6.483801e-08, 
    6.506309e-08, 6.510828e-08, 6.476632e-08, 6.497628e-08, 6.430245e-08, 
    6.441132e-08, 6.434649e-08, 6.410971e-08, 6.486627e-08, 6.447801e-08, 
    6.519495e-08, 6.498462e-08, 6.559846e-08, 6.529319e-08, 6.589279e-08, 
    6.614913e-08, 6.639036e-08, 6.667229e-08, 6.428748e-08, 6.420513e-08, 
    6.435257e-08, 6.455657e-08, 6.474583e-08, 6.499745e-08, 6.502319e-08, 
    6.507033e-08, 6.519242e-08, 6.529509e-08, 6.508524e-08, 6.532083e-08, 
    6.443658e-08, 6.489997e-08, 6.4174e-08, 6.439262e-08, 6.454454e-08, 
    6.44779e-08, 6.482399e-08, 6.490557e-08, 6.523705e-08, 6.506569e-08, 
    6.608587e-08, 6.563452e-08, 6.688694e-08, 6.653695e-08, 6.417636e-08, 
    6.428719e-08, 6.467292e-08, 6.448939e-08, 6.501424e-08, 6.514343e-08, 
    6.524845e-08, 6.538271e-08, 6.53972e-08, 6.547674e-08, 6.53464e-08, 
    6.547159e-08, 6.499798e-08, 6.520963e-08, 6.462883e-08, 6.47702e-08, 
    6.470516e-08, 6.463382e-08, 6.485399e-08, 6.508855e-08, 6.509355e-08, 
    6.516876e-08, 6.538072e-08, 6.501637e-08, 6.614414e-08, 6.544767e-08, 
    6.440805e-08, 6.462153e-08, 6.465201e-08, 6.456932e-08, 6.513049e-08, 
    6.492716e-08, 6.54748e-08, 6.532679e-08, 6.55693e-08, 6.544879e-08, 
    6.543107e-08, 6.527629e-08, 6.517993e-08, 6.493648e-08, 6.473839e-08, 
    6.458131e-08, 6.461784e-08, 6.479039e-08, 6.51029e-08, 6.539852e-08, 
    6.533376e-08, 6.555087e-08, 6.497619e-08, 6.521717e-08, 6.512403e-08, 
    6.536688e-08, 6.483475e-08, 6.528791e-08, 6.471893e-08, 6.476881e-08, 
    6.492312e-08, 6.523352e-08, 6.530218e-08, 6.537551e-08, 6.533025e-08, 
    6.511083e-08, 6.507487e-08, 6.491937e-08, 6.487644e-08, 6.475795e-08, 
    6.465985e-08, 6.474948e-08, 6.48436e-08, 6.511091e-08, 6.535181e-08, 
    6.561444e-08, 6.567871e-08, 6.598559e-08, 6.573579e-08, 6.614802e-08, 
    6.579756e-08, 6.640422e-08, 6.531416e-08, 6.578724e-08, 6.493014e-08, 
    6.502248e-08, 6.518949e-08, 6.557254e-08, 6.536574e-08, 6.560759e-08, 
    6.507346e-08, 6.479635e-08, 6.472464e-08, 6.459086e-08, 6.472769e-08, 
    6.471657e-08, 6.48475e-08, 6.480542e-08, 6.511979e-08, 6.495092e-08, 
    6.543063e-08, 6.560568e-08, 6.610003e-08, 6.640308e-08, 6.671156e-08, 
    6.684775e-08, 6.68892e-08, 6.690653e-08 ;

 SOILICE =
  57.57568, 57.76665, 57.72949, 57.88383, 57.79817, 57.8993, 57.61436, 
    57.77424, 57.67213, 57.59285, 58.18435, 57.89072, 58.49069, 58.30246, 
    58.77619, 58.46136, 58.83984, 58.7671, 58.98626, 58.92341, 59.20445, 
    59.01529, 59.35058, 59.15924, 59.18913, 59.00906, 57.94972, 58.14772, 
    57.938, 57.9662, 57.95354, 57.79994, 57.72265, 57.56111, 57.59041, 
    57.70908, 57.97888, 57.88718, 58.11854, 58.11331, 58.37177, 58.25512, 
    58.69092, 58.56682, 58.92603, 58.83552, 58.92178, 58.89561, 58.92212, 
    58.78942, 58.84624, 58.72959, 58.27695, 58.40969, 58.01453, 57.77799, 
    57.62136, 57.51043, 57.5261, 57.55598, 57.70977, 57.85469, 57.96534, 
    58.03945, 58.11256, 58.33429, 58.45195, 58.71603, 58.66832, 58.74918, 
    58.82652, 58.95656, 58.93514, 58.99249, 58.74705, 58.91007, 58.64115, 
    58.7146, 58.13242, 57.91191, 57.81837, 57.73663, 57.53815, 57.67515, 
    57.62111, 57.74975, 57.83162, 57.79112, 58.04148, 57.94403, 58.45893, 
    58.23668, 58.8175, 58.67811, 58.85095, 58.7627, 58.91397, 58.77782, 
    59.01384, 59.06534, 59.03014, 59.16544, 58.77028, 58.92177, 57.78999, 
    57.79659, 57.82736, 57.69218, 57.68393, 57.56031, 57.67029, 57.71718, 
    57.83637, 57.90697, 57.97414, 58.12208, 58.28767, 58.51988, 58.68714, 
    58.79946, 58.73056, 58.79139, 58.7234, 58.69156, 59.04604, 58.84677, 
    59.14597, 59.12938, 58.99385, 59.13124, 57.80122, 57.76323, 57.63147, 
    57.73456, 57.54686, 57.65186, 57.71231, 57.94606, 57.99754, 58.0453, 
    58.13972, 58.26109, 58.4745, 58.66067, 58.83102, 58.81853, 58.82293, 
    58.86103, 58.76668, 58.87654, 58.89499, 58.84675, 59.12716, 59.04694, 
    59.12902, 59.07678, 57.77558, 57.83953, 57.80497, 57.86998, 57.82417, 
    58.02811, 58.08938, 58.37678, 58.25869, 58.44673, 58.27777, 58.30768, 
    58.45286, 58.28689, 58.65039, 58.40375, 58.86251, 58.61554, 58.87802, 
    58.83029, 58.90934, 58.98021, 59.06947, 59.23446, 59.19622, 59.33441, 
    57.935, 58.01816, 58.01084, 58.09797, 58.16248, 58.30251, 58.52768, 
    58.44292, 58.59859, 58.62987, 58.39341, 58.53851, 58.07388, 58.14873, 
    58.10416, 57.94155, 58.46244, 58.19463, 58.6899, 58.54428, 58.9701, 
    58.75801, 59.17518, 59.35424, 59.52318, 59.72108, 58.06359, 58.00704, 
    58.10834, 58.24873, 58.37926, 58.55316, 58.57097, 58.60359, 58.68816, 
    58.75934, 58.61391, 58.77719, 58.1661, 58.48573, 57.98566, 58.13586, 
    58.24045, 58.19456, 58.43324, 58.48961, 58.71909, 58.60039, 59.31, 
    58.99518, 59.87214, 59.62601, 57.98729, 58.0634, 58.32895, 58.20248, 
    58.56479, 58.65421, 58.727, 58.82014, 58.83021, 58.88546, 58.79494, 
    58.88189, 58.55353, 58.70008, 58.29855, 58.39608, 58.3512, 58.30199, 
    58.45396, 58.61619, 58.61967, 58.67175, 58.81873, 58.56626, 59.35072, 
    58.86523, 58.1465, 58.2935, 58.31453, 58.25753, 58.64524, 58.50454, 
    58.88412, 58.78134, 58.94982, 58.86605, 58.85373, 58.7463, 58.6795, 
    58.51098, 58.37413, 58.2658, 58.29097, 58.41002, 58.62613, 58.83112, 
    58.78616, 58.937, 58.53845, 58.7053, 58.64077, 58.80916, 58.44067, 
    58.75433, 58.36069, 58.39513, 58.50174, 58.71663, 58.76426, 58.81514, 
    58.78374, 58.63162, 58.60673, 58.49915, 58.46947, 58.38763, 58.31994, 
    58.38178, 58.44678, 58.63169, 58.79869, 58.98122, 59.02596, 59.23993, 
    59.06569, 59.35344, 59.10872, 59.53286, 58.77255, 59.10154, 58.5066, 
    58.57048, 58.68612, 58.95206, 58.80836, 58.97644, 58.60576, 58.41413, 
    58.36464, 58.27238, 58.36675, 58.35907, 58.44948, 58.42041, 58.63783, 
    58.52098, 58.85342, 58.97512, 59.31992, 59.53209, 59.74871, 59.84454, 
    59.87373, 59.88594,
  78.79401, 79.09358, 79.03531, 79.27738, 79.14309, 79.30166, 78.85474, 
    79.10543, 78.94536, 78.82104, 79.74866, 79.28822, 80.2299, 79.93448, 
    80.67837, 80.18378, 80.77841, 80.66424, 81.00867, 80.90989, 81.35136, 
    81.05431, 81.58123, 81.28043, 81.32737, 81.04449, 79.38087, 79.69117, 
    79.36247, 79.40666, 79.38686, 79.14581, 79.02444, 78.77126, 78.8172, 
    79.00324, 79.42654, 79.28275, 79.64587, 79.63766, 80.04332, 79.86021, 
    80.54455, 80.34966, 80.91402, 80.77177, 80.9073, 80.8662, 80.90784, 
    80.6993, 80.78858, 80.60533, 79.89445, 80.10282, 79.48253, 79.11117, 
    78.86569, 78.69175, 78.71632, 78.76315, 79.00433, 79.23178, 79.40543, 
    79.52172, 79.63647, 79.98418, 80.16907, 80.58392, 80.50908, 80.63602, 
    80.75763, 80.96194, 80.92831, 81.01839, 80.63277, 80.88884, 80.46644, 
    80.58177, 79.66713, 79.32155, 79.17455, 79.04649, 78.73521, 78.95004, 
    78.86528, 79.06715, 79.19557, 79.13206, 79.5249, 79.37197, 80.18003, 
    79.83118, 80.74344, 80.52444, 80.79601, 80.65738, 80.895, 80.68112, 
    81.05199, 81.13286, 81.07758, 81.29028, 80.66927, 80.90724, 79.13026, 
    79.14061, 79.18892, 78.97674, 78.96381, 78.76997, 78.94248, 79.01599, 
    79.20307, 79.31379, 79.4192, 79.65137, 79.9112, 80.27582, 80.53862, 
    80.71513, 80.6069, 80.70244, 80.59562, 80.54562, 81.10251, 80.78938, 
    81.25967, 81.2336, 81.02052, 81.23654, 79.14789, 79.08831, 78.88157, 
    79.04333, 78.74889, 78.91352, 79.00827, 79.37504, 79.45595, 79.53085, 
    79.67908, 79.86957, 80.20457, 80.49699, 80.76473, 80.7451, 80.75201, 
    80.81185, 80.6636, 80.83621, 80.86516, 80.78941, 81.23011, 81.10402, 
    81.23305, 81.15095, 79.10769, 79.208, 79.15378, 79.25574, 79.18385, 
    79.50377, 79.59989, 80.05105, 79.86579, 80.16094, 79.89577, 79.94268, 
    80.17035, 79.91013, 80.48074, 80.09334, 80.81417, 80.42587, 80.83855, 
    80.76357, 80.88779, 80.99911, 81.13943, 81.39869, 81.33862, 81.55589, 
    79.3578, 79.48821, 79.47682, 79.61355, 79.71477, 79.93462, 80.28812, 
    80.15508, 80.39956, 80.44866, 80.07736, 80.30509, 79.57567, 79.69305, 
    79.62322, 79.36802, 80.18558, 79.76511, 80.54295, 80.31422, 80.98322, 
    80.64986, 81.30554, 81.58685, 81.85278, 82.16385, 79.55958, 79.47086, 
    79.62985, 79.85005, 80.05508, 80.32814, 80.35618, 80.40739, 80.54028, 
    80.65209, 80.42348, 80.68015, 79.72009, 80.22221, 79.43726, 79.67283, 
    79.8371, 79.76511, 80.13992, 80.22841, 80.58874, 80.40239, 81.51726, 
    81.02249, 82.40166, 82.01434, 79.43987, 79.55932, 79.97604, 79.77757, 
    80.34645, 80.48689, 80.6013, 80.74755, 80.76344, 80.85021, 80.70803, 
    80.84464, 80.32873, 80.55897, 79.92844, 80.0815, 80.01109, 79.93385, 
    80.17243, 80.42705, 80.43266, 80.5144, 80.7448, 80.34877, 81.58097, 
    80.81796, 79.68974, 79.9203, 79.95348, 79.86404, 80.47279, 80.2518, 
    80.84812, 80.68665, 80.95139, 80.81974, 80.80038, 80.63161, 80.52663, 
    80.26189, 80.04701, 79.87703, 79.91654, 80.10336, 80.44268, 80.76479, 
    80.69412, 80.93125, 80.30509, 80.5671, 80.46571, 80.73034, 80.15151, 
    80.6437, 80.02601, 80.08006, 80.24742, 80.58478, 80.65982, 80.73969, 
    80.69043, 80.45134, 80.41229, 80.24339, 80.19671, 80.0683, 79.96203, 
    80.05907, 80.16106, 80.45151, 80.71384, 81.00067, 81.07106, 81.40702, 
    81.13322, 81.58521, 81.20046, 81.86756, 80.67255, 81.1895, 80.2551, 
    80.35541, 80.53689, 80.95469, 80.7291, 80.99306, 80.41078, 80.10973, 
    80.03218, 79.88732, 80.0355, 80.02345, 80.16541, 80.11977, 80.46117, 
    80.27766, 80.79984, 80.99102, 81.53304, 81.86662, 82.20753, 82.3583, 
    82.40424, 82.42345,
  118.1172, 118.673, 118.5648, 119.0141, 118.7647, 119.0591, 118.2298, 
    118.695, 118.3979, 118.1672, 119.8895, 119.0342, 120.7661, 120.2339, 
    121.5725, 120.6833, 121.7525, 121.5469, 122.1666, 121.9888, 122.7838, 
    122.2487, 123.1976, 122.6559, 122.7405, 122.231, 119.206, 119.7828, 
    119.1719, 119.254, 119.2171, 118.7699, 118.5449, 118.0749, 118.1601, 
    118.5054, 119.2909, 119.0239, 119.6978, 119.6826, 120.4306, 120.0959, 
    121.3316, 120.981, 121.9962, 121.7403, 121.9842, 121.9102, 121.9851, 
    121.61, 121.7706, 121.4409, 120.1596, 120.5375, 119.3948, 118.7059, 
    118.2501, 117.9274, 117.973, 118.0599, 118.5074, 118.9293, 119.2515, 
    119.4674, 119.6804, 120.3248, 120.6567, 121.4025, 121.2677, 121.4962, 
    121.7149, 122.0825, 122.022, 122.1841, 121.4902, 121.9511, 121.191, 
    121.3985, 119.7382, 119.0959, 118.8235, 118.5856, 118.0081, 118.4066, 
    118.2494, 118.6238, 118.8621, 118.7442, 119.4733, 119.1894, 120.6764, 
    120.0422, 121.6893, 121.2954, 121.7839, 121.5345, 121.9621, 121.5772, 
    122.2446, 122.3902, 122.2907, 122.6735, 121.5559, 121.9841, 118.7409, 
    118.7601, 118.8497, 118.4562, 118.4322, 118.0725, 118.3925, 118.529, 
    118.8759, 119.0815, 119.2771, 119.7081, 120.1908, 120.8485, 121.3209, 
    121.6384, 121.4436, 121.6155, 121.4234, 121.3334, 122.3356, 121.7721, 
    122.6184, 122.5714, 122.188, 122.5767, 118.7736, 118.663, 118.2795, 
    118.5796, 118.0334, 118.3389, 118.5148, 119.1953, 119.3453, 119.4844, 
    119.7595, 120.1133, 120.7204, 121.2461, 121.7276, 121.6923, 121.7047, 
    121.8124, 121.5457, 121.8563, 121.9084, 121.772, 122.5652, 122.3382, 
    122.5704, 122.4226, 118.699, 118.8851, 118.7845, 118.9738, 118.8404, 
    119.4343, 119.6128, 120.4446, 120.1063, 120.642, 120.162, 120.2492, 
    120.6593, 120.1886, 121.217, 120.5207, 121.8166, 121.1185, 121.8605, 
    121.7255, 121.949, 122.1494, 122.4019, 122.8688, 122.7606, 123.1518, 
    119.1631, 119.4053, 119.384, 119.6379, 119.8259, 120.2341, 120.8705, 
    120.6313, 121.0707, 121.1591, 120.4916, 120.901, 119.5677, 119.7858, 
    119.6559, 119.1822, 120.6863, 119.9196, 121.3287, 120.9174, 122.1208, 
    121.5212, 122.701, 123.2079, 123.6865, 124.2474, 119.5377, 119.373, 
    119.6681, 120.0773, 120.4517, 120.9424, 120.9927, 121.0849, 121.3238, 
    121.525, 121.114, 121.5754, 119.8364, 120.7521, 119.3107, 119.7483, 
    120.0531, 119.9194, 120.604, 120.7631, 121.4112, 121.0758, 123.0826, 
    122.1917, 124.6758, 123.9779, 119.3154, 119.5372, 120.3097, 119.9425, 
    120.9752, 121.2279, 121.4335, 121.6968, 121.7253, 121.8815, 121.6256, 
    121.8714, 120.9434, 121.3575, 120.2225, 120.4991, 120.3725, 120.2326, 
    120.6625, 121.1204, 121.1303, 121.2774, 121.6927, 120.9794, 123.1979, 
    121.8242, 119.7793, 120.2078, 120.2691, 120.103, 121.2025, 120.8052, 
    121.8777, 121.5871, 122.0635, 121.8266, 121.7918, 121.4881, 121.2993, 
    120.8233, 120.4372, 120.1271, 120.2005, 120.5385, 121.1485, 121.7278, 
    121.6007, 122.0272, 120.9009, 121.3722, 121.1899, 121.6658, 120.6249, 
    121.5107, 120.3993, 120.4965, 120.7973, 121.4042, 121.5389, 121.6827, 
    121.5939, 121.164, 121.0937, 120.79, 120.7062, 120.4753, 120.2844, 
    120.4588, 120.6422, 121.1642, 121.6362, 122.1523, 122.2788, 122.8842, 
    122.3912, 123.2055, 122.5128, 123.7139, 121.5622, 122.4926, 120.811, 
    120.9913, 121.318, 122.0698, 121.6635, 122.1387, 121.091, 120.55, 
    120.4104, 120.1462, 120.4164, 120.3947, 120.6498, 120.5678, 121.1816, 
    120.8516, 121.7909, 122.135, 123.1108, 123.7117, 124.3258, 124.5976, 
    124.6804, 124.715,
  186.9664, 187.9677, 187.7727, 188.5826, 188.133, 188.6638, 187.1691, 
    188.0075, 187.4719, 187.0564, 190.1565, 188.6188, 191.7155, 190.757, 
    193.172, 191.5661, 193.4971, 193.1255, 194.2455, 193.9241, 195.3624, 
    194.394, 196.1112, 195.1308, 195.2839, 194.3621, 188.9286, 189.9695, 
    188.8671, 189.0152, 188.9487, 188.1423, 187.737, 186.89, 187.0435, 
    187.6657, 189.0818, 188.6001, 189.8158, 189.7883, 191.1098, 190.5161, 
    192.7365, 192.1033, 193.9375, 193.475, 193.9158, 193.782, 193.9175, 
    193.2395, 193.5298, 192.9339, 190.6272, 191.3029, 189.2691, 188.0273, 
    187.2058, 186.6246, 186.7066, 186.8632, 187.6693, 188.4296, 189.0106, 
    189.4, 189.7843, 190.9191, 191.5181, 192.8648, 192.6212, 193.034, 
    193.429, 194.0936, 193.9841, 194.2774, 193.0231, 193.856, 192.4825, 
    192.8574, 189.8891, 188.73, 188.2392, 187.8102, 186.7698, 187.4878, 
    187.2045, 187.879, 188.3085, 188.096, 189.4107, 188.8987, 191.5536, 
    190.4224, 193.3829, 192.6711, 193.5538, 193.103, 193.8759, 193.1802, 
    194.3866, 194.6501, 194.47, 195.1625, 193.1417, 193.9158, 188.09, 
    188.1247, 188.2862, 187.5771, 187.5338, 186.8858, 187.4623, 187.7082, 
    188.3334, 188.7041, 189.0569, 189.8344, 190.6818, 191.8642, 192.7172, 
    193.2907, 192.9389, 193.2495, 192.9023, 192.7397, 194.5514, 193.5325, 
    195.0628, 194.9778, 194.2844, 194.9874, 188.149, 187.9496, 187.2588, 
    187.7993, 186.8154, 187.3656, 187.6826, 188.9095, 189.1798, 189.4308, 
    189.9271, 190.5465, 191.6329, 192.5822, 193.452, 193.3881, 193.4106, 
    193.6053, 193.1233, 193.6845, 193.7789, 193.5323, 194.9665, 194.5559, 
    194.976, 194.7086, 188.0144, 188.3501, 188.1686, 188.5099, 188.2695, 
    189.3405, 189.6626, 191.1353, 190.5343, 191.4915, 190.6314, 190.7836, 
    191.5228, 190.6778, 192.5298, 191.2727, 193.6129, 192.352, 193.6921, 
    193.4482, 193.8522, 194.2146, 194.6712, 195.5161, 195.3201, 196.0283, 
    188.8512, 189.2882, 189.2496, 189.7076, 190.0451, 190.7572, 191.9039, 
    191.472, 192.2654, 192.425, 191.2199, 191.9591, 189.581, 189.9747, 
    189.7402, 188.8857, 191.5715, 190.2086, 192.7313, 191.9885, 194.1629, 
    193.0791, 195.2124, 196.1301, 196.9967, 198.0135, 189.5269, 189.2297, 
    189.7621, 190.4837, 191.1479, 192.0337, 192.1245, 192.2909, 192.7224, 
    193.0858, 192.3436, 193.177, 190.0637, 191.6902, 189.1174, 189.907, 
    190.4416, 190.2082, 191.4227, 191.7099, 192.8803, 192.2745, 195.9033, 
    194.2912, 198.7904, 197.5249, 189.1259, 189.5259, 190.8918, 190.2484, 
    192.093, 192.5492, 192.9207, 193.3964, 193.4478, 193.7302, 193.2676, 
    193.7119, 192.0356, 192.7833, 190.7371, 191.2335, 191.005, 190.7546, 
    191.5282, 192.3553, 192.3729, 192.6387, 193.3895, 192.1005, 196.1122, 
    193.627, 189.9628, 190.7115, 190.8184, 190.5284, 192.5034, 191.7859, 
    193.7233, 193.1982, 194.0592, 193.6309, 193.568, 193.0192, 192.6782, 
    191.8188, 191.1217, 190.5704, 190.6985, 191.3045, 192.4059, 193.4525, 
    193.2229, 193.9936, 191.9587, 192.81, 192.4806, 193.3403, 191.4606, 
    193.0605, 191.0533, 191.2286, 191.7717, 192.8678, 193.1109, 193.3709, 
    193.2104, 192.4339, 192.3069, 191.7585, 191.6073, 191.1904, 190.8459, 
    191.1607, 191.4917, 192.4342, 193.2868, 194.2197, 194.4486, 195.5443, 
    194.652, 196.1262, 194.8724, 197.0467, 193.1534, 194.8355, 191.7964, 
    192.122, 192.7121, 194.0707, 193.3362, 194.1954, 192.302, 191.3255, 
    191.0734, 190.6039, 191.0841, 191.045, 191.5054, 191.3574, 192.4656, 
    191.8697, 193.5664, 194.1886, 195.954, 197.0426, 198.1554, 198.6483, 
    198.7986, 198.8614,
  314.7132, 316.4507, 316.1121, 317.5188, 316.7377, 317.6599, 315.0646, 
    316.5199, 315.5901, 314.8691, 320.2661, 317.5817, 323.0769, 321.348, 
    325.708, 322.8074, 326.2959, 325.6238, 327.6396, 327.0685, 329.5956, 
    327.8995, 330.9085, 329.1897, 329.458, 327.8437, 318.12, 319.9308, 
    318.0131, 318.2706, 318.155, 316.7539, 316.0501, 314.5807, 314.8469, 
    315.9264, 318.3865, 317.5492, 319.663, 319.6151, 321.9841, 320.9139, 
    324.9208, 323.777, 327.0927, 326.2558, 327.0534, 326.8113, 327.0565, 
    325.83, 326.3549, 325.2776, 321.1141, 322.3324, 318.712, 316.5542, 
    315.1284, 314.1204, 314.2627, 314.5342, 315.9327, 317.2529, 318.2626, 
    318.9397, 319.6082, 321.6405, 322.7208, 325.1526, 324.7123, 325.4585, 
    326.1727, 327.3739, 327.177, 327.6954, 325.4387, 326.9452, 324.4618, 
    325.1392, 319.7908, 317.7749, 316.9222, 316.1772, 314.3722, 315.6176, 
    315.1261, 316.2966, 317.0426, 316.6734, 318.9583, 318.0681, 322.7849, 
    320.745, 326.0893, 324.8026, 326.3984, 325.5831, 326.9813, 325.7227, 
    327.8866, 328.3479, 328.0326, 329.2452, 325.6531, 327.0534, 316.6631, 
    316.7233, 317.0037, 315.7726, 315.6974, 314.5734, 315.5733, 316.0001, 
    317.0858, 317.7298, 318.3431, 319.6955, 321.2125, 323.3453, 324.8859, 
    325.9226, 325.2865, 325.848, 325.2204, 324.9266, 328.175, 326.3599, 
    329.0705, 328.9218, 327.7076, 328.9385, 316.7655, 316.4193, 315.2202, 
    316.1582, 314.4512, 315.4057, 315.9558, 318.0868, 318.5567, 318.9932, 
    319.8569, 320.9686, 322.9279, 324.6419, 326.2142, 326.0988, 326.1394, 
    326.4916, 325.6199, 326.635, 326.8057, 326.3596, 328.9018, 328.1829, 
    328.9186, 328.4503, 316.5318, 317.1147, 316.7996, 317.3925, 316.9747, 
    318.8364, 319.3965, 322.0302, 320.9467, 322.6727, 321.1216, 321.3959, 
    322.7294, 321.2052, 324.5473, 322.278, 326.5053, 324.2263, 326.6487, 
    326.2074, 326.9383, 327.5855, 328.3848, 329.8648, 329.5215, 330.763, 
    317.9856, 318.7453, 318.6782, 319.4749, 320.0652, 321.3484, 323.4169, 
    322.6375, 324.0696, 324.3579, 322.1826, 323.5166, 319.2546, 319.9396, 
    319.5315, 318.0455, 322.8171, 320.3598, 324.9114, 323.5696, 327.4951, 
    325.5401, 329.3326, 330.9417, 332.4626, 334.2497, 319.1605, 318.6435, 
    319.5697, 320.8556, 322.0528, 323.6514, 323.8153, 324.1158, 324.8953, 
    325.5521, 324.211, 325.717, 320.0989, 323.0312, 318.4483, 319.8218, 
    320.7796, 320.359, 322.5485, 323.0667, 325.1807, 324.0862, 330.5439, 
    327.7197, 335.6165, 333.3906, 318.4631, 319.1587, 321.5911, 320.4315, 
    323.7583, 324.5823, 325.2536, 326.1138, 326.2067, 326.7176, 325.8809, 
    326.6844, 323.6548, 325.0053, 321.312, 322.2073, 321.7951, 321.3437, 
    322.739, 324.2321, 324.2639, 324.7441, 326.1015, 323.7718, 330.9105, 
    326.5312, 319.9188, 321.2661, 321.4588, 320.9359, 324.4996, 323.204, 
    326.705, 325.7552, 327.3129, 326.538, 326.4241, 325.4317, 324.8154, 
    323.2633, 322.0057, 321.0117, 321.2426, 322.3354, 324.3236, 326.2152, 
    325.8, 327.1942, 323.516, 325.0535, 324.4585, 326.0122, 322.6169, 
    325.5066, 321.8823, 322.1984, 323.1783, 325.1582, 325.5975, 326.0676, 
    325.7774, 324.3741, 324.1447, 323.1544, 322.8816, 322.1296, 321.5083, 
    322.0759, 322.6731, 324.3747, 325.9156, 327.5946, 327.995, 329.9144, 
    328.3513, 330.9349, 328.7374, 332.5506, 325.6745, 328.6727, 323.2229, 
    323.8107, 324.8766, 327.3339, 326.0049, 327.552, 324.1357, 322.3732, 
    321.9185, 321.0721, 321.9379, 321.8673, 322.6978, 322.4307, 324.4313, 
    323.3552, 326.4213, 327.5401, 330.6327, 332.5432, 334.4991, 335.3664, 
    335.6308, 335.7415,
  523.2208, 526.4933, 525.8551, 528.509, 527.0347, 528.7755, 523.8821, 
    526.6239, 524.8715, 523.5142, 533.7062, 528.6277, 539.0436, 535.7582, 
    544.0582, 538.5309, 545.1812, 543.8974, 547.7717, 546.6583, 551.6522, 
    548.2866, 554.2629, 550.8459, 551.3788, 548.1761, 529.6447, 533.0709, 
    529.4426, 529.9293, 529.7108, 527.0652, 525.7383, 522.9714, 523.4724, 
    525.5051, 530.1483, 528.5663, 532.5637, 532.473, 536.966, 534.9344, 
    542.5559, 540.3761, 546.7047, 545.1046, 546.6295, 546.1664, 546.6355, 
    544.2911, 545.294, 543.2366, 535.3143, 537.6278, 530.7639, 526.6887, 
    524.0021, 522.1059, 522.3735, 522.884, 525.517, 528.0069, 529.9141, 
    531.1946, 532.4599, 536.3134, 538.3661, 542.9982, 542.1583, 543.5818, 
    544.9457, 547.2454, 546.866, 547.8823, 543.544, 546.4225, 541.6807, 
    542.9726, 532.8057, 528.9925, 527.3828, 525.9778, 522.5793, 524.9235, 
    523.9979, 526.2028, 527.6099, 526.9134, 531.2297, 529.5466, 538.4881, 
    534.6141, 544.7864, 542.3306, 545.377, 543.8198, 546.4915, 544.0862, 
    548.261, 549.1755, 548.5504, 550.9562, 543.9533, 546.6296, 526.8939, 
    527.0074, 527.5366, 525.2154, 525.0737, 522.9578, 524.84, 525.644, 
    527.6915, 528.9073, 530.0662, 532.6251, 535.501, 539.5542, 542.4893, 
    544.468, 543.2535, 544.3256, 543.1274, 542.5669, 548.8327, 545.3035, 
    550.6093, 550.314, 547.9066, 550.3473, 527.0872, 526.4342, 524.1751, 
    525.942, 522.728, 524.5242, 525.5605, 529.5819, 530.4702, 531.2958, 
    532.9308, 535.0382, 538.76, 542.0241, 545.0251, 544.8045, 544.8821, 
    545.5553, 543.89, 545.8293, 546.1557, 545.3029, 550.2745, 548.8483, 
    550.3077, 549.3785, 526.6463, 527.746, 527.1515, 528.2703, 527.4819, 
    530.999, 532.0591, 537.0537, 534.9967, 538.2747, 535.3284, 535.8491, 
    538.3826, 535.4871, 541.8438, 537.5245, 545.5815, 541.2319, 545.8555, 
    545.0121, 546.4093, 547.6646, 549.2487, 552.1871, 551.5048, 553.9733, 
    529.3906, 530.8268, 530.6999, 532.2073, 533.3256, 535.7589, 539.6904, 
    538.2078, 540.9333, 541.4827, 537.3432, 539.8803, 531.7904, 533.0875, 
    532.3146, 529.5039, 538.5493, 533.8839, 542.5381, 539.9812, 547.4854, 
    543.7376, 551.1298, 554.3289, 557.2599, 560.7106, 531.6123, 530.6342, 
    532.3868, 534.8238, 537.0966, 540.1368, 540.4489, 541.0213, 542.5072, 
    543.7606, 541.2027, 544.0753, 533.3893, 538.9565, 530.2653, 532.8645, 
    534.6797, 533.8823, 538.0386, 539.024, 543.0518, 540.9649, 553.5374, 
    547.9305, 563.3561, 559.0507, 530.2931, 531.6088, 536.2197, 534.0197, 
    540.3404, 541.9105, 543.1907, 544.8332, 545.0107, 545.9872, 544.3882, 
    545.9238, 540.1433, 542.717, 535.6899, 537.39, 536.607, 535.7499, 
    538.4006, 541.2429, 541.3035, 542.2189, 544.8098, 540.3661, 554.267, 
    545.6309, 533.0482, 535.6027, 535.9684, 534.9763, 541.7528, 539.2853, 
    545.9633, 544.1483, 547.126, 545.6438, 545.4262, 543.5308, 542.355, 
    539.3982, 537.007, 535.12, 535.558, 537.6334, 541.4173, 545.027, 
    544.2338, 546.899, 539.879, 542.8091, 541.6744, 544.6392, 538.1685, 
    543.6737, 536.7726, 537.3732, 539.2365, 543.0088, 543.8473, 544.7449, 
    544.1907, 541.5137, 541.0765, 539.191, 538.672, 537.2423, 536.0624, 
    537.1404, 538.2755, 541.5146, 544.4547, 547.6826, 548.476, 552.2856, 
    549.1824, 554.3157, 549.9484, 557.4296, 543.9943, 549.8199, 539.3213, 
    540.4402, 542.4717, 547.1663, 544.6252, 547.5983, 541.0593, 537.7054, 
    536.8413, 535.2346, 536.8781, 536.7442, 538.3223, 537.8145, 541.6226, 
    539.5729, 545.4208, 547.5746, 553.7141, 557.4154, 561.1931, 562.8717, 
    563.384, 563.5983,
  947.124, 953.9968, 952.6537, 958.2476, 955.1371, 958.8105, 948.5101, 
    954.2717, 950.5864, 947.7388, 969.1208, 958.4984, 980.1606, 973.3537, 
    990.6221, 979.096, 992.9768, 990.2852, 998.4262, 996.0811, 1006.634, 
    999.5121, 1012.188, 1004.924, 1006.054, 999.2789, 960.6486, 967.8129, 
    960.221, 961.2509, 960.7884, 955.2015, 952.4081, 946.6017, 947.6512, 
    951.9177, 961.7147, 958.3687, 966.7698, 966.5834, 975.8518, 971.6527, 
    987.4788, 982.932, 996.1787, 992.816, 996.0204, 995.0466, 996.0331, 
    991.1099, 993.2137, 988.9019, 972.4367, 977.2228, 963.019, 954.4083, 
    948.7616, 944.7905, 945.3502, 946.4188, 951.9427, 957.1875, 961.2188, 
    963.9323, 966.5566, 974.5015, 978.754, 988.4033, 986.6482, 989.6245, 
    992.4826, 997.3172, 996.5183, 998.6593, 989.5452, 995.5851, 985.6512, 
    988.3498, 967.2675, 959.2693, 955.8709, 952.9117, 945.7809, 950.6954, 
    948.7528, 953.3853, 956.3499, 954.8815, 964.0067, 960.4409, 979.0072, 
    970.9919, 992.1484, 987.0079, 993.3879, 990.1226, 995.7302, 990.6807, 
    999.4581, 1001.389, 1000.069, 1005.158, 990.4023, 996.0206, 954.8406, 
    955.0798, 956.1953, 951.3088, 951.0112, 946.5731, 950.5201, 952.2098, 
    956.522, 959.0893, 961.5409, 966.8961, 972.8223, 981.2219, 987.3397, 
    991.4807, 988.9374, 991.1822, 988.6735, 987.5017, 1000.665, 993.2335, 
    1004.423, 1003.798, 998.7104, 1003.868, 955.2477, 953.8723, 949.1246, 
    952.8365, 946.092, 949.8573, 952.0343, 960.5157, 962.3965, 964.147, 
    967.5247, 971.8668, 979.5717, 986.368, 992.6492, 992.1864, 992.3494, 
    993.7623, 990.2696, 994.3379, 995.024, 993.2323, 1003.714, 1000.698, 
    1003.784, 1001.818, 954.319, 956.6371, 955.3833, 957.7435, 956.0798, 
    963.5175, 965.7331, 976.0334, 971.7811, 978.5643, 972.466, 973.5416, 
    978.7881, 972.7936, 985.9915, 977.0087, 993.8173, 984.715, 994.393, 
    992.6219, 995.5572, 998.2003, 1001.544, 1007.77, 1006.322, 1011.571, 
    960.1111, 963.1523, 962.8834, 966.0375, 968.337, 973.3551, 981.5052, 
    978.4255, 984.0927, 985.238, 976.6331, 981.9001, 965.1812, 967.8472, 
    966.2579, 960.3507, 979.1342, 969.4866, 987.4415, 982.11, 997.8227, 
    989.9506, 1005.526, 1012.329, 1018.81, 1026.488, 964.8157, 962.7442, 
    966.4064, 971.4244, 976.1221, 982.4338, 983.0836, 984.2761, 987.377, 
    989.9986, 984.6542, 990.6578, 968.4683, 979.9798, 961.9623, 967.3884, 
    971.1271, 969.4833, 978.0745, 980.1201, 988.5153, 984.1585, 1010.642, 
    998.761, 1032.287, 1022.788, 962.0213, 964.8085, 974.3076, 969.7665, 
    982.8576, 986.1307, 988.806, 992.2466, 992.6191, 994.6697, 991.3137, 
    994.5366, 982.4473, 987.8155, 973.2126, 976.73, 975.1088, 973.3365, 
    978.8256, 984.738, 984.8643, 986.7748, 992.1975, 982.9113, 1012.197, 
    993.9212, 967.7662, 973.0325, 973.7881, 971.739, 985.8016, 980.6629, 
    994.6195, 990.8108, 997.0656, 993.9482, 993.4912, 989.5176, 987.0589, 
    980.8976, 975.9368, 972.0356, 972.9401, 977.2344, 985.1017, 992.6532, 
    990.9899, 996.5876, 981.8974, 988.008, 985.6381, 991.8398, 978.3441, 
    989.8168, 975.4514, 976.6952, 980.5614, 988.4255, 990.1802, 992.0616, 
    990.8997, 985.3028, 984.3911, 980.4669, 979.3889, 976.4241, 973.9824, 
    976.213, 978.5659, 985.3048, 991.4528, 998.2382, 999.9117, 1007.98, 
    1001.404, 1012.301, 1003.024, 1019.186, 990.4882, 1002.752, 980.7377, 
    983.0655, 987.3029, 997.1504, 991.8104, 998.0605, 984.3553, 977.3836, 
    975.5938, 972.2721, 975.6699, 975.3928, 978.6631, 977.6099, 985.53, 
    981.2609, 993.4799, 998.0106, 1011.018, 1019.154, 1027.565, 1031.236, 
    1032.348, 1032.813,
  1829.886, 1849.348, 1845.52, 1861.544, 1852.608, 1863.169, 1833.785, 
    1850.133, 1839.651, 1831.614, 1893.766, 1862.268, 1928.089, 1906.809, 
    1960.685, 1924.735, 1968.115, 1959.626, 1985.501, 1977.986, 2012.206, 
    1988.998, 2030.642, 2006.59, 2010.298, 1988.246, 1868.489, 1889.765, 
    1867.249, 1870.237, 1868.894, 1852.792, 1844.821, 1828.42, 1831.367, 
    1843.427, 1871.585, 1861.894, 1886.584, 1886.016, 1914.574, 1901.55, 
    1950.842, 1936.753, 1978.298, 1967.606, 1977.792, 1974.687, 1977.833, 
    1962.22, 1968.865, 1955.287, 1903.971, 1918.857, 1875.385, 1850.523, 
    1834.495, 1823.349, 1824.913, 1827.906, 1843.498, 1858.491, 1870.144, 
    1878.052, 1885.935, 1910.37, 1923.66, 1953.728, 1948.255, 1957.552, 
    1966.552, 1981.941, 1979.383, 1986.25, 1957.303, 1976.403, 1945.158, 
    1953.561, 1888.101, 1864.494, 1854.71, 1846.254, 1826.119, 1839.96, 
    1834.47, 1847.603, 1856.084, 1851.876, 1878.27, 1867.887, 1924.456, 
    1899.514, 1965.496, 1949.374, 1969.418, 1959.115, 1976.866, 1960.869, 
    1988.823, 1995.068, 1990.795, 2007.355, 1959.994, 1977.793, 1851.759, 
    1852.443, 1855.64, 1841.698, 1840.854, 1828.339, 1839.463, 1844.257, 
    1856.578, 1863.974, 1871.08, 1886.969, 1905.163, 1931.441, 1950.408, 
    1963.389, 1955.399, 1962.448, 1954.573, 1950.913, 1992.722, 1968.928, 
    2004.948, 2002.904, 1986.415, 2003.134, 1852.924, 1848.992, 1835.518, 
    1846.04, 1826.99, 1837.588, 1843.758, 1868.104, 1873.57, 1878.68, 
    1888.885, 1902.211, 1926.232, 1947.383, 1967.079, 1965.616, 1966.13, 
    1970.605, 1959.577, 1972.432, 1974.615, 1968.924, 2002.631, 1992.829, 
    2002.861, 1996.46, 1850.268, 1856.909, 1853.312, 1860.092, 1855.309, 
    1876.84, 1883.43, 1915.14, 1901.946, 1923.064, 1904.061, 1907.391, 
    1923.767, 1905.074, 1946.214, 1918.187, 1970.779, 1942.257, 1972.608, 
    1966.992, 1976.314, 1984.775, 1995.569, 2015.952, 2011.177, 2028.578, 
    1866.931, 1875.773, 1874.989, 1884.355, 1891.367, 1906.813, 1932.338, 
    1922.628, 1940.333, 1943.876, 1917.013, 1933.58, 1881.755, 1889.87, 
    1885.026, 1867.625, 1924.855, 1894.888, 1950.725, 1934.225, 1983.562, 
    1958.575, 2008.563, 2031.113, 2053.028, 2079.233, 1880.647, 1874.583, 
    1885.478, 1900.846, 1915.417, 1935.22, 1937.22, 1940.9, 1950.524, 
    1958.726, 1942.069, 1960.797, 1891.769, 1927.518, 1872.306, 1888.469, 
    1899.93, 1894.877, 1921.526, 1927.961, 1954.078, 1940.536, 2025.48, 
    1986.578, 2099.502, 2066.699, 1872.477, 1880.625, 1909.768, 1895.746, 
    1936.524, 1946.646, 1954.987, 1965.806, 1966.983, 1973.487, 1962.862, 
    1973.064, 1935.261, 1951.892, 1906.371, 1917.316, 1912.259, 1906.755, 
    1923.885, 1942.328, 1942.719, 1948.649, 1965.651, 1936.689, 2030.671, 
    1971.109, 1889.622, 1905.814, 1908.155, 1901.816, 1945.624, 1929.674, 
    1973.328, 1961.279, 1981.135, 1971.195, 1969.745, 1957.216, 1949.533, 
    1930.416, 1914.839, 1902.732, 1905.528, 1918.894, 1943.454, 1967.091, 
    1961.842, 1979.605, 1933.571, 1952.493, 1945.117, 1964.521, 1922.372, 
    1958.155, 1913.326, 1917.207, 1929.354, 1953.797, 1959.296, 1965.221, 
    1961.558, 1944.077, 1941.255, 1929.055, 1925.657, 1916.36, 1908.758, 
    1915.701, 1923.069, 1944.083, 1963.301, 1984.896, 1990.287, 2016.643, 
    1995.115, 2031.019, 2000.38, 2054.315, 1960.264, 1999.495, 1929.911, 
    1937.164, 1950.293, 1981.406, 1964.428, 1984.326, 1941.145, 1919.361, 
    1913.769, 1903.462, 1914.007, 1913.143, 1923.374, 1920.069, 1944.782, 
    1931.565, 1969.709, 1984.165, 2026.734, 2054.207, 2082.894, 2095.755, 
    2099.718, 2101.382,
  5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597,
  8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILLIQ =
  4.547437, 4.565955, 4.56235, 4.577317, 4.56901, 4.578816, 4.551187, 
    4.566692, 4.556789, 4.549101, 4.606462, 4.577985, 4.636159, 4.617906, 
    4.663849, 4.633317, 4.670022, 4.662964, 4.684221, 4.678125, 4.705389, 
    4.687037, 4.719559, 4.701001, 4.703902, 4.686432, 4.583704, 4.602911, 
    4.582568, 4.585303, 4.584075, 4.569182, 4.561691, 4.546023, 4.548864, 
    4.560372, 4.586533, 4.57764, 4.600072, 4.599565, 4.624626, 4.613315, 
    4.655575, 4.643537, 4.678379, 4.669601, 4.677967, 4.675429, 4.678, 
    4.66513, 4.670641, 4.659326, 4.615432, 4.628304, 4.589988, 4.567058, 
    4.551866, 4.541109, 4.542628, 4.545527, 4.56044, 4.57449, 4.585217, 
    4.592403, 4.599492, 4.620997, 4.632403, 4.658013, 4.653382, 4.661228, 
    4.668728, 4.681341, 4.679263, 4.684826, 4.661019, 4.676833, 4.650746, 
    4.657872, 4.601428, 4.580037, 4.570973, 4.563043, 4.543797, 4.557083, 
    4.551842, 4.564314, 4.572253, 4.568325, 4.5926, 4.583152, 4.63308, 
    4.611529, 4.667853, 4.654333, 4.671097, 4.662537, 4.677211, 4.664003, 
    4.686897, 4.691893, 4.688479, 4.701601, 4.663272, 4.677968, 4.568215, 
    4.568856, 4.571839, 4.558734, 4.557933, 4.545945, 4.55661, 4.561158, 
    4.572712, 4.579558, 4.586072, 4.600416, 4.616473, 4.638988, 4.655208, 
    4.666102, 4.65942, 4.665319, 4.658725, 4.655636, 4.690021, 4.670693, 
    4.699712, 4.698102, 4.684959, 4.698284, 4.569305, 4.565621, 4.552846, 
    4.562841, 4.544641, 4.554823, 4.560686, 4.583352, 4.58834, 4.592971, 
    4.602126, 4.613894, 4.634587, 4.652642, 4.669164, 4.667952, 4.668379, 
    4.672076, 4.662923, 4.673579, 4.67537, 4.67069, 4.697887, 4.690106, 
    4.698069, 4.693001, 4.566818, 4.57302, 4.569668, 4.575973, 4.571531, 
    4.591308, 4.597248, 4.625114, 4.613662, 4.631895, 4.615511, 4.618412, 
    4.632494, 4.616395, 4.651647, 4.62773, 4.672219, 4.648268, 4.673723, 
    4.669093, 4.67676, 4.683635, 4.692292, 4.708296, 4.704587, 4.71799, 
    4.582276, 4.590341, 4.589629, 4.598078, 4.604333, 4.617909, 4.639742, 
    4.631524, 4.646618, 4.649653, 4.626723, 4.640794, 4.595743, 4.603003, 
    4.598678, 4.582913, 4.633419, 4.607452, 4.655477, 4.641352, 4.682655, 
    4.662085, 4.702546, 4.719917, 4.736298, 4.755495, 4.594745, 4.589261, 
    4.599082, 4.612699, 4.625352, 4.642213, 4.64394, 4.647104, 4.655307, 
    4.662211, 4.648107, 4.663943, 4.604691, 4.635677, 4.58719, 4.601756, 
    4.611894, 4.607443, 4.630585, 4.636051, 4.658309, 4.646792, 4.715627, 
    4.68509, 4.770141, 4.746274, 4.587346, 4.594726, 4.620475, 4.608211, 
    4.64334, 4.652015, 4.659074, 4.66811, 4.669086, 4.674446, 4.665664, 
    4.674098, 4.642249, 4.656464, 4.617525, 4.626983, 4.62263, 4.617859, 
    4.632594, 4.648329, 4.648663, 4.653717, 4.667983, 4.643482, 4.719583, 
    4.672492, 4.602782, 4.61704, 4.619076, 4.613548, 4.651145, 4.637498, 
    4.674314, 4.664345, 4.680687, 4.672562, 4.671367, 4.660946, 4.654467, 
    4.638124, 4.624855, 4.614349, 4.61679, 4.628335, 4.649292, 4.669175, 
    4.664815, 4.679443, 4.640786, 4.656971, 4.650712, 4.667044, 4.631306, 
    4.661735, 4.62355, 4.626889, 4.637228, 4.658072, 4.662688, 4.667625, 
    4.664578, 4.649825, 4.647409, 4.636976, 4.634099, 4.626162, 4.619599, 
    4.625596, 4.631899, 4.64983, 4.666029, 4.683733, 4.688072, 4.708832, 
    4.691931, 4.719847, 4.696112, 4.737245, 4.663498, 4.69541, 4.637698, 
    4.643892, 4.655111, 4.680908, 4.666967, 4.683272, 4.647315, 4.628735, 
    4.623933, 4.614988, 4.624138, 4.623393, 4.632159, 4.629341, 4.650426, 
    4.639091, 4.671338, 4.683143, 4.716585, 4.737165, 4.75817, 4.767464, 
    4.770294, 4.771478,
  5.63329, 5.656574, 5.652041, 5.670864, 5.660416, 5.67275, 5.638004, 
    5.657501, 5.645048, 5.635382, 5.707526, 5.671704, 5.744902, 5.721928, 
    5.779763, 5.741323, 5.787535, 5.778648, 5.805419, 5.79774, 5.832085, 
    5.808966, 5.849941, 5.826556, 5.830211, 5.808205, 5.678897, 5.703058, 
    5.677469, 5.680909, 5.679364, 5.660632, 5.651212, 5.631512, 5.635084, 
    5.649554, 5.682456, 5.671269, 5.699488, 5.698849, 5.730386, 5.716151, 
    5.769344, 5.754189, 5.798061, 5.787005, 5.797542, 5.794345, 5.797584, 
    5.781375, 5.788316, 5.774067, 5.718815, 5.735014, 5.686802, 5.657961, 
    5.638858, 5.625334, 5.627244, 5.630888, 5.649639, 5.667308, 5.680801, 
    5.689841, 5.698758, 5.725818, 5.740173, 5.772414, 5.766583, 5.776462, 
    5.785906, 5.801791, 5.799174, 5.806181, 5.776199, 5.796113, 5.763265, 
    5.772236, 5.701193, 5.674285, 5.662885, 5.652913, 5.628714, 5.645417, 
    5.638828, 5.654511, 5.664495, 5.659555, 5.690088, 5.678204, 5.741024, 
    5.713903, 5.784804, 5.76778, 5.788889, 5.778111, 5.796589, 5.779956, 
    5.80879, 5.815083, 5.810782, 5.827312, 5.779036, 5.797543, 5.659417, 
    5.660223, 5.663975, 5.647494, 5.646486, 5.631414, 5.644823, 5.650541, 
    5.665073, 5.673683, 5.681876, 5.699921, 5.720125, 5.748462, 5.768882, 
    5.7826, 5.774185, 5.781614, 5.77331, 5.769421, 5.812725, 5.788381, 
    5.824933, 5.822906, 5.806348, 5.823134, 5.660788, 5.656154, 5.64009, 
    5.652658, 5.629775, 5.642577, 5.649948, 5.678453, 5.684729, 5.690555, 
    5.702072, 5.716879, 5.742922, 5.765651, 5.786456, 5.784929, 5.785467, 
    5.790122, 5.778597, 5.792016, 5.794271, 5.788377, 5.822634, 5.812832, 
    5.822862, 5.816479, 5.65766, 5.66546, 5.661244, 5.669173, 5.663587, 
    5.688462, 5.695935, 5.730999, 5.716588, 5.739534, 5.718915, 5.722565, 
    5.740288, 5.720027, 5.764398, 5.734292, 5.790303, 5.760145, 5.792197, 
    5.786366, 5.796021, 5.804681, 5.815586, 5.835748, 5.831075, 5.847963, 
    5.677101, 5.687246, 5.68635, 5.696979, 5.704849, 5.721932, 5.749412, 
    5.739067, 5.758068, 5.761888, 5.733024, 5.750735, 5.694041, 5.703175, 
    5.697734, 5.677902, 5.741452, 5.708774, 5.76922, 5.751438, 5.803446, 
    5.777541, 5.828503, 5.850392, 5.871037, 5.895238, 5.692786, 5.685887, 
    5.698243, 5.715375, 5.731299, 5.752522, 5.754696, 5.75868, 5.769006, 
    5.7777, 5.759942, 5.779881, 5.705298, 5.744294, 5.683282, 5.701606, 
    5.714363, 5.708763, 5.737885, 5.744765, 5.772786, 5.758287, 5.844985, 
    5.806513, 5.913707, 5.883612, 5.683478, 5.692762, 5.725161, 5.709728, 
    5.75394, 5.764862, 5.773749, 5.785128, 5.786356, 5.793107, 5.782048, 
    5.792669, 5.752567, 5.770463, 5.721449, 5.733352, 5.727873, 5.721869, 
    5.740414, 5.760221, 5.760642, 5.767005, 5.784967, 5.754119, 5.84997, 
    5.790646, 5.702898, 5.720838, 5.723401, 5.716444, 5.763766, 5.746587, 
    5.792942, 5.780386, 5.800967, 5.790734, 5.78923, 5.776107, 5.767949, 
    5.747375, 5.730673, 5.717453, 5.720524, 5.735054, 5.761434, 5.786469, 
    5.780979, 5.799401, 5.750726, 5.771102, 5.763221, 5.783785, 5.738792, 
    5.777099, 5.729032, 5.733234, 5.746246, 5.772488, 5.778301, 5.784517, 
    5.78068, 5.762104, 5.759064, 5.745929, 5.742308, 5.732318, 5.724059, 
    5.731606, 5.73954, 5.762111, 5.782508, 5.804804, 5.810269, 5.836423, 
    5.81513, 5.850302, 5.820396, 5.872231, 5.77932, 5.819512, 5.746838, 
    5.754635, 5.76876, 5.801246, 5.783689, 5.804224, 5.758944, 5.735557, 
    5.729513, 5.718256, 5.729771, 5.728834, 5.739866, 5.736319, 5.762861, 
    5.748593, 5.789193, 5.80406, 5.846193, 5.87213, 5.898612, 5.91033, 
    5.9139, 5.915393,
  8.097958, 8.132158, 8.1255, 8.153154, 8.137803, 8.155926, 8.10488, 8.13352, 
    8.115227, 8.101029, 8.207046, 8.154389, 8.262018, 8.228224, 8.313323, 
    8.256754, 8.324766, 8.311683, 8.351101, 8.339793, 8.390382, 8.356324, 
    8.416696, 8.382236, 8.387621, 8.355203, 8.164961, 8.200477, 8.162861, 
    8.167916, 8.165647, 8.138121, 8.124281, 8.095345, 8.100592, 8.121845, 
    8.170191, 8.153751, 8.195228, 8.194289, 8.240664, 8.219728, 8.297988, 
    8.275683, 8.340264, 8.323986, 8.3395, 8.334793, 8.339561, 8.315697, 
    8.325915, 8.304939, 8.223646, 8.247472, 8.176579, 8.134196, 8.106135, 
    8.086273, 8.089079, 8.09443, 8.12197, 8.147929, 8.167759, 8.181046, 
    8.194154, 8.233946, 8.255061, 8.302505, 8.293924, 8.308463, 8.322368, 
    8.345758, 8.341904, 8.352222, 8.308077, 8.337397, 8.28904, 8.302244, 
    8.197734, 8.158183, 8.14143, 8.12678, 8.091237, 8.115769, 8.106091, 
    8.129128, 8.143796, 8.136539, 8.181409, 8.163941, 8.256314, 8.216423, 
    8.320745, 8.295685, 8.32676, 8.31089, 8.338098, 8.313608, 8.356065, 
    8.365335, 8.358999, 8.38335, 8.312253, 8.339501, 8.136335, 8.137519, 
    8.143032, 8.118819, 8.11734, 8.095202, 8.114897, 8.123296, 8.144646, 
    8.157297, 8.169338, 8.195864, 8.225573, 8.267257, 8.297307, 8.3175, 
    8.305113, 8.316049, 8.303824, 8.2981, 8.361861, 8.326012, 8.379845, 
    8.376858, 8.352468, 8.377194, 8.13835, 8.131541, 8.107945, 8.126407, 
    8.092794, 8.111596, 8.122425, 8.164309, 8.173532, 8.182095, 8.199026, 
    8.220798, 8.259107, 8.292552, 8.323176, 8.32093, 8.32172, 8.328575, 
    8.311606, 8.331363, 8.334683, 8.326005, 8.376458, 8.36202, 8.376794, 
    8.367391, 8.133754, 8.145214, 8.13902, 8.150671, 8.142462, 8.179018, 
    8.190004, 8.241567, 8.22037, 8.254122, 8.223793, 8.229161, 8.25523, 
    8.225429, 8.290708, 8.24641, 8.328841, 8.284448, 8.33163, 8.323044, 
    8.337262, 8.350014, 8.366076, 8.39578, 8.388893, 8.413781, 8.162321, 
    8.177232, 8.175916, 8.191539, 8.20311, 8.22823, 8.268655, 8.253434, 
    8.281391, 8.287013, 8.244545, 8.270601, 8.187221, 8.200648, 8.19265, 
    8.163498, 8.256943, 8.20888, 8.297805, 8.271636, 8.348194, 8.310053, 
    8.385105, 8.41736, 8.447794, 8.483485, 8.185375, 8.175234, 8.193398, 
    8.218587, 8.242007, 8.273231, 8.276429, 8.282291, 8.29749, 8.310287, 
    8.284148, 8.313497, 8.20377, 8.261124, 8.171405, 8.198341, 8.217099, 
    8.208863, 8.251695, 8.261817, 8.303052, 8.281714, 8.409392, 8.352713, 
    8.510731, 8.466338, 8.171694, 8.18534, 8.232979, 8.210284, 8.275317, 
    8.291389, 8.304471, 8.321222, 8.32303, 8.33297, 8.316688, 8.332325, 
    8.273297, 8.299633, 8.22752, 8.245027, 8.236968, 8.228138, 8.255415, 
    8.28456, 8.28518, 8.294544, 8.320984, 8.275581, 8.416738, 8.329345, 
    8.200241, 8.226622, 8.23039, 8.22016, 8.289777, 8.264498, 8.332726, 
    8.314241, 8.344544, 8.329475, 8.327261, 8.307942, 8.295934, 8.265656, 
    8.241086, 8.221642, 8.22616, 8.24753, 8.286345, 8.323195, 8.315113, 
    8.342238, 8.270588, 8.300574, 8.288976, 8.319245, 8.253031, 8.309402, 
    8.238672, 8.244854, 8.263997, 8.302614, 8.311171, 8.320323, 8.314674, 
    8.287332, 8.282857, 8.26353, 8.258203, 8.243507, 8.231359, 8.242458, 
    8.254129, 8.287341, 8.317365, 8.350196, 8.358244, 8.396774, 8.365404, 
    8.417227, 8.37316, 8.449554, 8.312672, 8.371859, 8.264868, 8.27634, 
    8.297128, 8.344954, 8.319102, 8.34934, 8.282681, 8.24827, 8.239381, 
    8.222824, 8.239759, 8.23838, 8.25461, 8.249393, 8.288445, 8.267449, 
    8.327207, 8.3491, 8.411171, 8.449406, 8.488461, 8.50575, 8.511017, 8.51322,
  12.66457, 12.72004, 12.70924, 12.7541, 12.72919, 12.7586, 12.6758, 
    12.72225, 12.69257, 12.66955, 12.84161, 12.75611, 12.93096, 12.87602, 
    13.01443, 12.9224, 13.03306, 13.01176, 13.07595, 13.05753, 13.13997, 
    13.08446, 13.18289, 13.12669, 13.13547, 13.08264, 12.77326, 12.83093, 
    12.76986, 12.77806, 12.77438, 12.72971, 12.70726, 12.66034, 12.66884, 
    12.70331, 12.78175, 12.75507, 12.82241, 12.82088, 12.89624, 12.86221, 
    12.98947, 12.95318, 13.0583, 13.03179, 13.05706, 13.04939, 13.05716, 
    13.0183, 13.03493, 13.00079, 12.86858, 12.9073, 12.79213, 12.72334, 
    12.67783, 12.64563, 12.65018, 12.65886, 12.70351, 12.74562, 12.77781, 
    12.79938, 12.82067, 12.88531, 12.91964, 12.99682, 12.98286, 13.00652, 
    13.02916, 13.06725, 13.06097, 13.07778, 13.00589, 13.05363, 12.97491, 
    12.9964, 12.82648, 12.76226, 12.73508, 12.71131, 12.65368, 12.69345, 
    12.67776, 12.71512, 12.73892, 12.72714, 12.79997, 12.77161, 12.92168, 
    12.85684, 13.02652, 12.98572, 13.03631, 13.01047, 13.05477, 13.0149, 
    13.08404, 13.09914, 13.08882, 13.12851, 13.01269, 13.05706, 12.72681, 
    12.72873, 12.73768, 12.6984, 12.696, 12.66011, 12.69204, 12.70566, 
    12.7403, 12.76083, 12.78037, 12.82344, 12.87171, 12.93948, 12.98837, 
    13.02123, 13.00107, 13.01887, 12.99897, 12.98965, 13.09348, 13.03509, 
    13.12279, 13.11793, 13.07818, 13.11847, 12.73008, 12.71904, 12.68077, 
    12.71071, 12.6562, 12.68669, 12.70425, 12.77221, 12.78718, 12.80108, 
    12.82858, 12.86395, 12.92622, 12.98063, 13.03047, 13.02682, 13.0281, 
    13.03926, 13.01164, 13.0438, 13.04921, 13.03508, 13.11727, 13.09374, 
    13.11782, 13.1025, 12.72262, 12.74122, 12.73117, 12.75007, 12.73675, 
    12.79609, 12.81393, 12.8977, 12.86325, 12.91812, 12.86882, 12.87754, 
    12.91992, 12.87147, 12.97762, 12.90558, 13.0397, 12.96744, 13.04424, 
    13.03026, 13.05341, 13.07418, 13.10035, 13.14877, 13.13754, 13.17813, 
    12.76898, 12.79319, 12.79105, 12.81642, 12.83521, 12.87603, 12.94175, 
    12.917, 12.96247, 12.97161, 12.90255, 12.94492, 12.80941, 12.83121, 
    12.81822, 12.77089, 12.9227, 12.84459, 12.98917, 12.9466, 13.07122, 
    13.00911, 13.13137, 13.18397, 13.23363, 13.29191, 12.80641, 12.78994, 
    12.81944, 12.86036, 12.89842, 12.94919, 12.9544, 12.96393, 12.98866, 
    13.00949, 12.96695, 13.01472, 12.83628, 12.9295, 12.78373, 12.82747, 
    12.85794, 12.84456, 12.91417, 12.93063, 12.99771, 12.96299, 13.17097, 
    13.07858, 13.33643, 13.26391, 12.78419, 12.80635, 12.88375, 12.84687, 
    12.95259, 12.97873, 13.00002, 13.02729, 13.03024, 13.04642, 13.01991, 
    13.04537, 12.9493, 12.99215, 12.87487, 12.90333, 12.89023, 12.87588, 
    12.92022, 12.96762, 12.96863, 12.98387, 13.0269, 12.95302, 13.18295, 
    13.04052, 12.83055, 12.87341, 12.87954, 12.86291, 12.97611, 12.93499, 
    13.04603, 13.01593, 13.06527, 13.04073, 13.03712, 13.00567, 12.98613, 
    12.93687, 12.89692, 12.86532, 12.87266, 12.9074, 12.97053, 13.03051, 
    13.01735, 13.06152, 12.94489, 12.99368, 12.97481, 13.02407, 12.91634, 
    13.00805, 12.893, 12.90305, 12.93417, 12.997, 13.01093, 13.02583, 
    13.01663, 12.97213, 12.96485, 12.93342, 12.92475, 12.90086, 12.88111, 
    12.89915, 12.91813, 12.97215, 13.02101, 13.07448, 13.08759, 13.15039, 
    13.09926, 13.18375, 13.1119, 13.2365, 13.01337, 13.10978, 12.93559, 
    12.95425, 12.98807, 13.06594, 13.02384, 13.07308, 12.96457, 12.9086, 
    12.89415, 12.86724, 12.89477, 12.89252, 12.91891, 12.91043, 12.97394, 
    12.93979, 13.03704, 13.07269, 13.17387, 13.23626, 13.30004, 13.32829, 
    13.3369, 13.3405,
  20.59555, 20.6916, 20.67289, 20.75065, 20.70747, 20.75845, 20.61498, 
    20.69543, 20.64403, 20.60417, 20.90253, 20.75413, 21.05791, 20.96234, 
    21.20336, 21.04301, 21.23585, 21.1987, 21.31072, 21.27856, 21.4226, 
    21.32558, 21.49769, 21.39938, 21.41473, 21.32239, 20.78389, 20.88399, 
    20.77798, 20.79221, 20.78582, 20.70836, 20.66946, 20.58822, 20.60294, 
    20.66262, 20.79862, 20.75233, 20.86919, 20.86654, 20.9975, 20.93834, 
    21.15984, 21.09661, 21.2799, 21.23364, 21.27773, 21.26435, 21.2779, 
    21.2101, 21.23912, 21.17956, 20.9494, 21.01675, 20.81661, 20.69733, 
    20.6185, 20.56278, 20.57064, 20.58566, 20.66297, 20.73595, 20.79177, 
    20.8292, 20.86616, 20.9785, 21.03822, 21.17266, 21.14831, 21.18956, 
    21.22904, 21.29552, 21.28456, 21.31391, 21.18847, 21.27175, 21.13446, 
    21.17191, 20.87625, 20.7648, 20.71767, 20.67648, 20.5767, 20.64555, 
    20.61838, 20.68308, 20.72432, 20.70391, 20.83022, 20.78102, 21.04177, 
    20.929, 21.22443, 21.15331, 21.24152, 21.19645, 21.27374, 21.20417, 
    21.32484, 21.35123, 21.3332, 21.40255, 21.20032, 21.27773, 20.70334, 
    20.70667, 20.72218, 20.65412, 20.64996, 20.58782, 20.6431, 20.66669, 
    20.72671, 20.76231, 20.79622, 20.87098, 20.95484, 21.07274, 21.15791, 
    21.21522, 21.18005, 21.21109, 21.1764, 21.16016, 21.34134, 21.23939, 
    21.39256, 21.38405, 21.31461, 21.38501, 20.70901, 20.68987, 20.62358, 
    20.67544, 20.58107, 20.63383, 20.66425, 20.78205, 20.80803, 20.83216, 
    20.8799, 20.94136, 21.04967, 21.14442, 21.23134, 21.22495, 21.2272, 
    21.24667, 21.19848, 21.2546, 21.26403, 21.23937, 21.38291, 21.34179, 
    21.38387, 21.35708, 20.69608, 20.72831, 20.71089, 20.74366, 20.72057, 
    20.82349, 20.85446, 21.00005, 20.94015, 21.03556, 20.94982, 20.96498, 
    21.0387, 20.95444, 21.13919, 21.01375, 21.24743, 21.12144, 21.25536, 
    21.23096, 21.27136, 21.30763, 21.35334, 21.43799, 21.41836, 21.48936, 
    20.77645, 20.81845, 20.81474, 20.85878, 20.89142, 20.96235, 21.0767, 
    21.03362, 21.11278, 21.12872, 21.00847, 21.08222, 20.84661, 20.88448, 
    20.86192, 20.77977, 21.04355, 20.90771, 21.15932, 21.08515, 21.30245, 
    21.19407, 21.40756, 21.49958, 21.58658, 21.68879, 20.84141, 20.81282, 
    20.86403, 20.93511, 21.0013, 21.08966, 21.09872, 21.11534, 21.15843, 
    21.19474, 21.1206, 21.20385, 20.89328, 21.05538, 20.80204, 20.87797, 
    20.93091, 20.90766, 21.0287, 21.05734, 21.17421, 21.1137, 21.47684, 
    21.3153, 21.76696, 21.63965, 20.80285, 20.8413, 20.97577, 20.91167, 
    21.09557, 21.14113, 21.17823, 21.22579, 21.23092, 21.25916, 21.21291, 
    21.25733, 21.08985, 21.16451, 20.96035, 21.00983, 20.98705, 20.96209, 
    21.03922, 21.12177, 21.12352, 21.15007, 21.22511, 21.09632, 21.4978, 
    21.24886, 20.88333, 20.95781, 20.96846, 20.93955, 21.13655, 21.06493, 
    21.25847, 21.20597, 21.29207, 21.24924, 21.24294, 21.18808, 21.15401, 
    21.06821, 20.99869, 20.94374, 20.9565, 21.01692, 21.12682, 21.23139, 
    21.20844, 21.28551, 21.08218, 21.16718, 21.13428, 21.22017, 21.03248, 
    21.19222, 20.99187, 21.00935, 21.06351, 21.17296, 21.19725, 21.22323, 
    21.20719, 21.12962, 21.11694, 21.06219, 21.04711, 21.00554, 20.9712, 
    21.00257, 21.03559, 21.12965, 21.21483, 21.30815, 21.33105, 21.44083, 
    21.35143, 21.4992, 21.37352, 21.59161, 21.20151, 21.36981, 21.06598, 
    21.09847, 21.1574, 21.29324, 21.21977, 21.30571, 21.11644, 21.01901, 
    20.99387, 20.94708, 20.99494, 20.99104, 21.03695, 21.02218, 21.13278, 
    21.07329, 21.24279, 21.30503, 21.48191, 21.59119, 21.70305, 21.75266, 
    21.76778, 21.77411,
  34.63898, 34.81974, 34.78448, 34.93107, 34.84964, 34.94579, 34.67551, 
    34.82695, 34.73016, 34.65519, 35.21814, 34.93763, 35.51294, 35.33147, 
    35.78992, 35.48462, 35.85194, 35.78104, 35.99503, 35.93353, 36.20937, 
    36.02347, 36.35357, 36.16483, 36.19426, 36.01736, 34.9938, 35.18304, 
    34.98264, 35.00952, 34.99745, 34.85132, 34.77803, 34.62521, 34.65288, 
    34.76515, 35.02161, 34.93423, 35.15502, 35.15001, 35.39818, 35.28597, 
    35.70694, 35.58654, 35.93609, 35.84771, 35.93194, 35.90636, 35.93227, 
    35.80278, 35.85817, 35.74453, 35.30695, 35.43474, 35.05562, 34.83053, 
    34.68213, 34.5774, 34.59218, 34.62038, 34.76581, 34.90334, 35.00868, 
    35.07941, 35.1493, 35.36214, 35.47552, 35.73137, 35.68498, 35.7636, 
    35.83894, 35.96596, 35.945, 36.00114, 35.76151, 35.92051, 35.6586, 
    35.72995, 35.1684, 34.95778, 34.86886, 34.79126, 34.60355, 34.73302, 
    34.6819, 34.80369, 34.88141, 34.84294, 35.08134, 34.98838, 35.48226, 
    35.26828, 35.83014, 35.69449, 35.86276, 35.77674, 35.92432, 35.79146, 
    36.02205, 36.07257, 36.03804, 36.17092, 35.78412, 35.93194, 34.84186, 
    34.84813, 34.87736, 34.74915, 34.74133, 34.62445, 34.72841, 34.77283, 
    34.88592, 34.95307, 35.01708, 35.15842, 35.31726, 35.54114, 35.70326, 
    35.81255, 35.74547, 35.80468, 35.7385, 35.70755, 36.05363, 35.8587, 
    36.15176, 36.13545, 36.00248, 36.13729, 34.85254, 34.81647, 34.69169, 
    34.78928, 34.61176, 34.71098, 34.76822, 34.99033, 35.03939, 35.085, 
    35.1753, 35.2917, 35.49728, 35.67757, 35.84332, 35.83113, 35.83543, 
    35.8726, 35.78062, 35.88774, 35.90577, 35.85867, 36.13327, 36.05449, 
    36.1351, 36.08378, 34.82819, 34.88893, 34.85609, 34.91788, 34.87434, 
    35.0686, 35.12716, 35.40303, 35.28941, 35.47047, 35.30774, 35.33649, 
    35.47643, 35.3165, 35.6676, 35.42903, 35.87405, 35.6338, 35.88919, 
    35.8426, 35.91978, 35.98911, 36.07661, 36.23891, 36.20123, 36.33757, 
    34.97977, 35.05909, 35.05208, 35.13534, 35.19711, 35.33151, 35.54867, 
    35.46677, 35.61732, 35.64766, 35.41902, 35.55915, 35.11231, 35.18396, 
    35.14127, 34.98602, 35.48564, 35.22794, 35.70595, 35.56473, 35.97921, 
    35.77221, 36.18051, 36.35721, 36.52464, 36.72184, 35.10248, 35.04845, 
    35.14526, 35.27986, 35.4054, 35.57332, 35.59056, 35.62218, 35.70425, 
    35.77348, 35.63219, 35.79086, 35.20063, 35.50813, 35.02807, 35.17164, 
    35.2719, 35.22786, 35.45743, 35.51186, 35.73433, 35.61906, 36.31349, 
    36.0038, 36.87302, 36.62698, 35.02961, 35.10229, 35.35696, 35.23545, 
    35.58456, 35.67129, 35.742, 35.83272, 35.84253, 35.89646, 35.80815, 
    35.89296, 35.57368, 35.71584, 35.3277, 35.4216, 35.37835, 35.33101, 
    35.47742, 35.63441, 35.63776, 35.68833, 35.83143, 35.58599, 36.35379, 
    35.87679, 35.18179, 35.32288, 35.34308, 35.28828, 35.66258, 35.52629, 
    35.89514, 35.79489, 35.95936, 35.87749, 35.86547, 35.76078, 35.69584, 
    35.53252, 35.40045, 35.29622, 35.32042, 35.43505, 35.64405, 35.84343, 
    35.79961, 35.94682, 35.55908, 35.72092, 35.65825, 35.82201, 35.4646, 
    35.76868, 35.3875, 35.42068, 35.52359, 35.73195, 35.77826, 35.82785, 
    35.79724, 35.64937, 35.62523, 35.52108, 35.49241, 35.41345, 35.34827, 
    35.40782, 35.47051, 35.64943, 35.81181, 35.9901, 36.03392, 36.24435, 
    36.07294, 36.35648, 36.11526, 36.53433, 35.78639, 36.10815, 35.52828, 
    35.59008, 35.70229, 35.96159, 35.82123, 35.98545, 35.62428, 35.43902, 
    35.3913, 35.30255, 35.39333, 35.38593, 35.4731, 35.44505, 35.65539, 
    35.54218, 35.86518, 35.98414, 36.32325, 36.53352, 36.7494, 36.84534, 
    36.87461, 36.88686,
  60.67812, 61.07083, 60.99409, 61.31372, 61.13599, 61.34589, 60.75732, 
    61.08654, 60.87596, 60.71325, 61.9436, 61.32805, 62.59598, 62.19373, 
    63.21417, 62.53307, 63.35332, 63.19427, 63.67535, 63.53676, 64.1604, 
    63.73952, 64.48857, 64.05934, 64.12612, 63.72573, 61.45091, 61.86631, 
    61.42648, 61.48533, 61.4589, 61.13967, 60.98005, 60.64828, 60.70824, 
    60.95203, 61.51183, 61.32064, 61.80466, 61.79365, 62.34135, 62.09321, 
    63.02843, 62.75974, 63.54253, 63.34382, 63.53318, 63.47564, 63.53393, 
    63.243, 63.36732, 63.11252, 62.13955, 62.42237, 61.58636, 61.09434, 
    60.77169, 60.54478, 60.57676, 60.63782, 60.95346, 61.25315, 61.48349, 
    61.63854, 61.79207, 62.26156, 62.51286, 63.08306, 62.97935, 63.15522, 
    63.32412, 63.60981, 63.5626, 63.68912, 63.15054, 63.50746, 62.92043, 
    63.0799, 61.83408, 61.3721, 61.17791, 61.00883, 60.60137, 60.88219, 
    60.77119, 61.03589, 61.20528, 61.12138, 61.6428, 61.43905, 62.52781, 
    62.05416, 63.30437, 63.0006, 63.37762, 63.18466, 63.51603, 63.21764, 
    63.73633, 63.85044, 63.77242, 64.07315, 63.20119, 63.5332, 61.11904, 
    61.13271, 61.19645, 60.91724, 60.90023, 60.64664, 60.87217, 60.96872, 
    61.21512, 61.36182, 61.5019, 61.81213, 62.16233, 62.65869, 63.02021, 
    63.26492, 63.11462, 63.24727, 63.09903, 63.02979, 63.80764, 63.36849, 
    64.02972, 63.99276, 63.69214, 63.99692, 61.14231, 61.06372, 60.79243, 
    61.00454, 60.61915, 60.8343, 60.95869, 61.44333, 61.55079, 61.65081, 
    61.84928, 62.10587, 62.56117, 62.96279, 63.33397, 63.30662, 63.31625, 
    63.39974, 63.19335, 63.43375, 63.4743, 63.36842, 63.98781, 63.80959, 
    63.99197, 63.8758, 61.08924, 61.22169, 61.15005, 61.28492, 61.18986, 
    61.61485, 61.7434, 62.35209, 62.1008, 62.50164, 62.14127, 62.20483, 
    62.51487, 62.16063, 62.94054, 62.40972, 63.40299, 62.86511, 63.43701, 
    63.33235, 63.50581, 63.66199, 63.85958, 64.22751, 64.14191, 64.4521, 
    61.4202, 61.59398, 61.57861, 61.76139, 61.89728, 62.19381, 62.67543, 
    62.49344, 62.82833, 62.89602, 62.38752, 62.69877, 61.71079, 61.86834, 
    61.77442, 61.43389, 62.53532, 61.96521, 63.02622, 62.71117, 63.63968, 
    63.17449, 64.09491, 64.49689, 64.87986, 65.33361, 61.68919, 61.57066, 
    61.7832, 62.07972, 62.35733, 62.7303, 62.7687, 62.83917, 63.02241, 
    63.17733, 62.86152, 63.21629, 61.90504, 62.58529, 61.52598, 61.84122, 
    62.06215, 61.96502, 62.4727, 62.59358, 63.08968, 62.83222, 64.39722, 
    63.69513, 65.68346, 65.11497, 61.52935, 61.68877, 62.2501, 61.98175, 
    62.75535, 62.94876, 63.10686, 63.31018, 63.33219, 63.45336, 63.25504, 
    63.44549, 62.7311, 63.04832, 62.18539, 62.39325, 62.29745, 62.19272, 
    62.51709, 62.86647, 62.87393, 62.98683, 63.30727, 62.75852, 64.48909, 
    63.40913, 61.86355, 62.17475, 62.2194, 62.09832, 62.92932, 62.62566, 
    63.4504, 63.22533, 63.59494, 63.41073, 63.38372, 63.14891, 63.00362, 
    62.63952, 62.34638, 62.11584, 62.16929, 62.42306, 62.88795, 63.3342, 
    63.23591, 63.5667, 62.69861, 63.0597, 62.91965, 63.28613, 62.48863, 
    63.16659, 62.31769, 62.39119, 62.61966, 63.08437, 63.18806, 63.29924, 
    63.23058, 62.89984, 62.84597, 62.61407, 62.55037, 62.37517, 62.23088, 
    62.3627, 62.50174, 62.89996, 63.26327, 63.66423, 63.76313, 64.23988, 
    63.8513, 64.49522, 63.94703, 64.90211, 63.20626, 63.93095, 62.63008, 
    62.76763, 63.01803, 63.59995, 63.2844, 63.65374, 62.84386, 62.43187, 
    62.3261, 62.12982, 62.33061, 62.31422, 62.50748, 62.44524, 62.91327, 
    62.66099, 63.38306, 63.65079, 64.41946, 64.90024, 65.39728, 65.61928, 
    65.68716, 65.71558,
  116.3177, 117.5456, 117.3041, 118.3151, 117.7513, 118.4176, 116.5637, 
    117.5951, 116.9338, 116.4267, 120.3481, 118.3608, 122.5137, 121.171, 
    124.6257, 122.3021, 125.1096, 124.5568, 126.2417, 125.7524, 127.9808, 
    126.4694, 129.1813, 127.615, 127.8565, 126.4205, 118.7533, 120.0957, 
    118.6751, 118.8636, 118.7789, 117.7629, 117.26, 116.2252, 116.4112, 
    117.1721, 118.9486, 118.3372, 119.895, 119.8591, 121.6609, 120.8392, 
    123.9848, 123.0673, 125.7727, 125.0765, 125.7398, 125.5376, 125.7424, 
    124.7257, 125.1585, 124.2743, 120.992, 121.9312, 119.1884, 117.6198, 
    116.6085, 115.9052, 116.004, 116.1928, 117.1766, 118.1225, 118.8577, 
    119.3567, 119.854, 121.3957, 122.2342, 124.1727, 123.8163, 124.4217, 
    125.0078, 126.0099, 125.8434, 126.2906, 124.4055, 125.6493, 123.6146, 
    124.1618, 119.9907, 118.5013, 117.8839, 117.3504, 116.08, 116.9533, 
    116.6069, 117.4356, 117.9706, 117.7051, 119.3704, 118.7153, 122.2844, 
    120.7108, 124.939, 123.8892, 125.1944, 124.5235, 125.6795, 124.6378, 
    126.4581, 126.8647, 126.5865, 127.6649, 124.5807, 125.7398, 117.6977, 
    117.7409, 117.9426, 117.063, 117.0098, 116.2201, 116.922, 117.2244, 
    118.0018, 118.4685, 118.9168, 119.9193, 121.0672, 122.7252, 123.9565, 
    124.8018, 124.2815, 124.7406, 124.2277, 123.9894, 126.712, 125.1625, 
    127.5082, 127.375, 126.3013, 127.39, 117.7713, 117.5232, 116.6731, 
    117.3369, 116.135, 116.8037, 117.193, 118.729, 119.0739, 119.3963, 
    120.0402, 120.8809, 122.3965, 123.7596, 125.0421, 124.9468, 124.9804, 
    125.2717, 124.5536, 125.3907, 125.5329, 125.1623, 127.3572, 126.7189, 
    127.3722, 126.9554, 117.6037, 118.0227, 117.7958, 118.2235, 117.9217, 
    119.2802, 119.696, 121.6967, 120.8642, 122.1966, 120.9977, 121.2077, 
    122.241, 121.0616, 123.6834, 121.8889, 125.2831, 123.4257, 125.4021, 
    125.0365, 125.6435, 126.1945, 126.8974, 128.2247, 127.9137, 129.0469, 
    118.655, 119.2129, 119.1634, 119.7544, 120.1967, 121.1713, 122.7818, 
    122.1691, 123.3005, 123.5312, 121.8148, 122.8607, 119.5903, 120.1023, 
    119.7967, 118.6988, 122.3096, 120.4189, 123.9772, 122.9027, 126.1155, 
    124.4883, 127.7435, 129.212, 130.6391, 132.3671, 119.5204, 119.1378, 
    119.8252, 120.7948, 121.7141, 122.9675, 123.0977, 123.3373, 123.9641, 
    124.4982, 123.4135, 124.6331, 120.2221, 122.4777, 118.9941, 120.0139, 
    120.737, 120.4182, 122.0996, 122.5056, 124.1955, 123.3137, 128.8451, 
    126.3119, 133.7281, 131.5293, 119.0049, 119.519, 121.3577, 120.4731, 
    123.0524, 123.7116, 124.2547, 124.9592, 125.0359, 125.4594, 124.7675, 
    125.4319, 122.9702, 124.0532, 121.1434, 121.8339, 121.5149, 121.1676, 
    122.2484, 123.4304, 123.4558, 123.842, 124.9491, 123.0632, 129.1832, 
    125.3046, 120.0867, 121.1082, 121.256, 120.856, 123.645, 122.6137, 
    125.4491, 124.6644, 125.9574, 125.3102, 125.2157, 124.3999, 123.8996, 
    122.6605, 121.6777, 120.9138, 121.0902, 121.9335, 123.5037, 125.0429, 
    124.7011, 125.8578, 122.8601, 124.0923, 123.612, 124.8756, 122.153, 
    124.461, 121.5822, 121.8271, 122.5935, 124.1772, 124.5353, 124.9212, 
    124.6826, 123.5443, 123.3605, 122.5746, 122.3602, 121.7736, 121.294, 
    121.7321, 122.1969, 123.5447, 124.7961, 126.2024, 126.5534, 128.2697, 
    126.8678, 129.2058, 127.2107, 130.7228, 124.5983, 127.153, 122.6286, 
    123.0941, 123.9491, 125.9751, 124.8695, 126.1652, 123.3533, 121.963, 
    121.6102, 120.9599, 121.6252, 121.5707, 122.2162, 122.0077, 123.5901, 
    122.733, 125.2134, 126.1548, 128.9268, 130.7158, 132.6128, 133.4764, 
    133.7426, 133.8543,
  366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466,
  603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILPSI =
  -0.02010258, -0.01977483, -0.0198381, -0.01957703, -0.01972141, 
    -0.01955111, -0.02003568, -0.01976193, -0.01993623, -0.02007286, 
    -0.01908082, -0.01956547, -0.01859121, -0.01889026, -0.01814875, 
    -0.01863739, -0.01805192, -0.01816269, -0.01783159, -0.01792577, 
    -0.01750933, -0.0177883, -0.01729765, -0.01757554, -0.01753174, 
    -0.01779758, -0.01946692, -0.01914043, -0.01948644, -0.01943947, 
    -0.01946054, -0.0197184, -0.01984971, -0.02012789, -0.02007709, 
    -0.01987294, -0.01941839, -0.01957145, -0.01918825, -0.01919682, 
    -0.01877947, -0.01896642, -0.01827957, -0.01847202, -0.01792183, 
    -0.0180585, -0.01792822, -0.01796762, -0.01792771, -0.01812861, 
    -0.01804224, -0.01822013, -0.01893124, -0.01871918, -0.01935933, 
    -0.01975552, -0.02002358, -0.02021614, -0.0201888, -0.02013678, 
    -0.01987175, -0.01962602, -0.01944094, -0.01931818, -0.01919805, 
    -0.01883919, -0.01865227, -0.01824091, -0.01831445, -0.01819008, 
    -0.01807217, -0.01787601, -0.01790814, -0.01782228, -0.01819337, 
    -0.01794581, -0.01835647, -0.01824315, -0.01916539, -0.01953004, 
    -0.01968716, -0.01982592, -0.0201678, -0.01993103, -0.020024, -0.0198036, 
    -0.01966489, -0.01973336, -0.01931483, -0.0194764, -0.01864126, 
    -0.01899615, -0.01808587, -0.01829933, -0.01803512, -0.01816943, 
    -0.01793995, -0.01814633, -0.01779045, -0.01771395, -0.01776619, 
    -0.01756647, -0.01815785, -0.01792821, -0.01973528, -0.01972409, 
    -0.01967208, -0.01990183, -0.01991599, -0.02012928, -0.01993939, 
    -0.0198591, -0.01965689, -0.0195383, -0.01942629, -0.01918245, 
    -0.01891399, -0.0185454, -0.01828541, -0.01811333, -0.01821865, 
    -0.01812563, -0.01822964, -0.01827862, -0.01774256, -0.01804143, 
    -0.01759505, -0.01761943, -0.01782024, -0.01761668, -0.01971624, 
    -0.01978069, -0.02000615, -0.01982947, -0.02015266, -0.01997104, 
    -0.01986741, -0.01947298, -0.01938748, -0.01930853, -0.01915364, 
    -0.0189568, -0.01861674, -0.01832624, -0.01806534, -0.01808432, 
    -0.01807763, -0.01801984, -0.01816334, -0.0179964, -0.01796854, 
    -0.01804148, -0.0176227, -0.01774126, -0.01761995, -0.01769704, 
    -0.01975972, -0.01965154, -0.01970991, -0.01960029, -0.01967744, 
    -0.01933684, -0.01923597, -0.01877145, -0.01896064, -0.01866054, 
    -0.01892993, -0.01888189, -0.01865078, -0.01891528, -0.0183421, 
    -0.01872857, -0.0180176, -0.01839609, -0.01799416, -0.01806645, 
    -0.01794694, -0.01784062, -0.01770785, -0.01746564, -0.01752141, 
    -0.01732094, -0.01949147, -0.01935332, -0.01936546, -0.01922194, 
    -0.01911652, -0.0188902, -0.01853321, -0.0186666, -0.01842253, 
    -0.01837394, -0.01874507, -0.01851623, -0.01926147, -0.01913888, 
    -0.01921178, -0.01948052, -0.01863573, -0.01906422, -0.01828114, 
    -0.01850722, -0.01785574, -0.01817655, -0.01755219, -0.01729235, 
    -0.01705171, -0.01677497, -0.01927839, -0.01937175, -0.01920495, 
    -0.01897667, -0.01876755, -0.01849334, -0.01846554, -0.01841473, 
    -0.01828384, -0.01817456, -0.01839867, -0.01814728, -0.01911052, 
    -0.01859905, -0.01940715, -0.01915987, -0.01899006, -0.01906437, 
    -0.01868192, -0.01859298, -0.01823623, -0.01841973, -0.01735607, 
    -0.01781822, -0.01656761, -0.0169072, -0.01940448, -0.01927872, 
    -0.01884781, -0.01905153, -0.0184752, -0.01833624, -0.01822412, 
    -0.01808184, -0.01806657, -0.01798292, -0.01812021, -0.01798833, 
    -0.01849276, -0.01826548, -0.01889656, -0.01874081, -0.0188123, 
    -0.01889103, -0.01864916, -0.01839512, -0.01838977, -0.01830912, 
    -0.01808384, -0.01847291, -0.0172973, -0.01801335, -0.01914259, 
    -0.01890459, -0.01887091, -0.01896254, -0.01835012, -0.01856951, 
    -0.01798496, -0.01814096, -0.01788612, -0.01801226, -0.0180309, 
    -0.01819452, -0.01829719, -0.01855938, -0.01877572, -0.01894922, 
    -0.01890873, -0.01871867, -0.01837971, -0.01806517, -0.01813356, 
    -0.01790535, -0.01851635, -0.01825742, -0.01835702, -0.01809856, 
    -0.01867015, -0.01818208, -0.01879715, -0.01874234, -0.01857389, 
    -0.01823998, -0.01816704, -0.01808944, -0.01813729, -0.0183712, 
    -0.01840984, -0.01857798, -0.01862467, -0.01875426, -0.01886227, 
    -0.01876355, -0.01866047, -0.01837111, -0.01811448, -0.01783911, 
    -0.01777242, -0.0174576, -0.01771337, -0.0172934, -0.01764967, 
    -0.01703792, -0.01815428, -0.01766035, -0.01856628, -0.01846632, 
    -0.01828695, -0.0178827, -0.01809976, -0.01784621, -0.01841136, 
    -0.01871213, -0.01879086, -0.01893862, -0.01878749, -0.01879974, 
    -0.01865624, -0.01870223, -0.01836159, -0.01854373, -0.01803136, 
    -0.01784821, -0.01734182, -0.01703908, -0.01673686, -0.01660528, 
    -0.01656546, -0.01654884,
  -0.05392879, -0.05288604, -0.0530871, -0.05225819, -0.05271635, 
    -0.05217599, -0.05371569, -0.05284504, -0.05339914, -0.0538341, 
    -0.05068813, -0.05222154, -0.04914599, -0.05008706, -0.04775852, 
    -0.04929113, -0.04745567, -0.04780213, -0.04676764, -0.04706157, 
    -0.04576404, -0.04663264, -0.04510658, -0.04596996, -0.04583371, 
    -0.04666157, -0.05190917, -0.05087638, -0.05197102, -0.05182223, 
    -0.05188896, -0.0527068, -0.05312401, -0.05400945, -0.05384757, 
    -0.05319784, -0.05175547, -0.05224048, -0.05102742, -0.05105449, 
    -0.04973809, -0.05032713, -0.04816814, -0.04877164, -0.04704926, 
    -0.04747625, -0.04706921, -0.04719226, -0.0470676, -0.04769551, 
    -0.0474254, -0.04798193, -0.05021623, -0.04954835, -0.05156849, 
    -0.05282469, -0.05367717, -0.05429079, -0.0542036, -0.05403776, 
    -0.05319406, -0.05241357, -0.05182686, -0.05143826, -0.05105838, 
    -0.04992617, -0.04933792, -0.04804701, -0.0482774, -0.04788786, 
    -0.04751896, -0.04690623, -0.04700652, -0.0467386, -0.04789817, 
    -0.04712413, -0.04840914, -0.04805402, -0.05095523, -0.05210918, 
    -0.05260764, -0.05304838, -0.05413665, -0.0533826, -0.05367852, 
    -0.05297742, -0.05253691, -0.05275431, -0.05142767, -0.05193919, 
    -0.04930329, -0.05042091, -0.04756183, -0.04823003, -0.04740315, 
    -0.04782321, -0.04710582, -0.04775095, -0.04663933, -0.04640089, 
    -0.04656368, -0.04594174, -0.04778698, -0.04706917, -0.0527604, 
    -0.05272487, -0.05255973, -0.05328974, -0.05333477, -0.05401387, 
    -0.0534092, -0.05315384, -0.05251152, -0.05213538, -0.05178047, 
    -0.05100908, -0.05016184, -0.04900206, -0.04818641, -0.04764771, 
    -0.0479773, -0.04768619, -0.04801172, -0.04816513, -0.04649006, 
    -0.04742287, -0.04603065, -0.04610655, -0.04673224, -0.046098, 
    -0.05269995, -0.05290463, -0.05362168, -0.05305966, -0.05408838, 
    -0.05350994, -0.05318026, -0.05192836, -0.05165759, -0.05140772, 
    -0.05091806, -0.0502968, -0.04922621, -0.04831436, -0.0474976, 
    -0.04755696, -0.04753605, -0.04735541, -0.04780416, -0.04728216, 
    -0.04719511, -0.04742302, -0.04611673, -0.04648599, -0.04610817, 
    -0.04634821, -0.05283801, -0.05249456, -0.05267985, -0.05233197, 
    -0.05257677, -0.05149732, -0.05117825, -0.04971287, -0.05030893, 
    -0.04936392, -0.0502121, -0.05006067, -0.04933325, -0.0501659, 
    -0.0483641, -0.0495779, -0.0473484, -0.04853339, -0.04727516, 
    -0.04750111, -0.04712767, -0.04679581, -0.0463819, -0.04562822, 
    -0.04580159, -0.04517883, -0.05198694, -0.05154944, -0.05158788, 
    -0.05113389, -0.05080083, -0.05008687, -0.04896375, -0.04938296, 
    -0.04861632, -0.04846391, -0.04962982, -0.04891044, -0.05125887, 
    -0.05087145, -0.0511018, -0.05195225, -0.04928592, -0.05063571, 
    -0.04817304, -0.04888215, -0.04684297, -0.04784552, -0.04589732, 
    -0.04509013, -0.04434449, -0.04348934, -0.05131239, -0.05160779, 
    -0.0510802, -0.05035949, -0.04970058, -0.04883857, -0.04875131, 
    -0.04859186, -0.04818151, -0.04783929, -0.0485415, -0.04775392, 
    -0.05078189, -0.0491706, -0.05171987, -0.05093776, -0.0504017, 
    -0.05063619, -0.04943113, -0.04915152, -0.04803238, -0.04860755, 
    -0.04528788, -0.04672594, -0.04285018, -0.04389763, -0.05171141, 
    -0.05131344, -0.0499533, -0.05059566, -0.04878163, -0.0483457, 
    -0.04799443, -0.04754922, -0.04750146, -0.04724003, -0.04766923, 
    -0.04725693, -0.04883675, -0.04812397, -0.05010691, -0.04961641, 
    -0.04984145, -0.05008948, -0.04932813, -0.04853034, -0.04851355, 
    -0.04826071, -0.0475555, -0.04877442, -0.04510553, -0.04733514, 
    -0.05088316, -0.05013224, -0.05002608, -0.0503149, -0.04838922, 
    -0.04907779, -0.0472464, -0.04773413, -0.04693778, -0.04733172, 
    -0.04738997, -0.04790176, -0.04822332, -0.04904597, -0.04972629, 
    -0.05027292, -0.05014525, -0.04954675, -0.04848201, -0.04749709, 
    -0.047711, -0.04699781, -0.04891081, -0.04809874, -0.04841087, 
    -0.04760149, -0.04939412, -0.04786285, -0.04979375, -0.04962122, 
    -0.04909156, -0.04804411, -0.04781575, -0.04757299, -0.04772265, 
    -0.04845532, -0.04857653, -0.04910439, -0.04925114, -0.04965874, 
    -0.04999884, -0.04968798, -0.0493637, -0.04845505, -0.04765129, 
    -0.04679109, -0.04658313, -0.04560323, -0.04639909, -0.04509341, 
    -0.04620073, -0.04430184, -0.04777583, -0.04623395, -0.04906764, 
    -0.04875374, -0.04819123, -0.04692712, -0.04760527, -0.04681325, 
    -0.0485813, -0.04952618, -0.04977395, -0.05023948, -0.04976336, 
    -0.0498019, -0.04935039, -0.04949502, -0.04842519, -0.04899679, 
    -0.0473914, -0.04681948, -0.04524364, -0.04430543, -0.04337175, 
    -0.04296617, -0.04284354, -0.04279238,
  -0.07870831, -0.07705726, -0.07737544, -0.07606426, -0.0767888, 
    -0.07593434, -0.07837072, -0.0769924, -0.0778694, -0.07855829, 
    -0.07358485, -0.07600633, -0.07115486, -0.07263708, -0.06897327, 
    -0.07138334, -0.06849768, -0.06904177, -0.06741803, -0.06787911, 
    -0.06584527, -0.06720632, -0.06481629, -0.06616777, -0.06595436, 
    -0.0672517, -0.07551263, -0.07388186, -0.07561037, -0.07537525, 
    -0.0754807, -0.0767737, -0.07743385, -0.07883612, -0.07857963, 
    -0.07755072, -0.07526978, -0.07603627, -0.07412019, -0.0741629, 
    -0.0720872, -0.07301552, -0.06961685, -0.0705658, -0.06785981, 
    -0.06852999, -0.06789111, -0.0680842, -0.0678886, -0.06887429, 
    -0.06845015, -0.06932423, -0.07284068, -0.07178835, -0.07497443, 
    -0.07696021, -0.0783097, -0.07928204, -0.07914381, -0.07888098, 
    -0.07754473, -0.07630993, -0.07538258, -0.07476875, -0.07416904, 
    -0.07238355, -0.071457, -0.06942651, -0.0697886, -0.06917644, 
    -0.06859704, -0.06763541, -0.06779274, -0.06737249, -0.06919263, 
    -0.06797729, -0.0699957, -0.06943751, -0.07400628, -0.07582872, 
    -0.07661686, -0.07731415, -0.0790377, -0.07784322, -0.07831183, 
    -0.07720187, -0.07650498, -0.07684885, -0.07475204, -0.07556006, 
    -0.07140247, -0.0731634, -0.06866436, -0.06971414, -0.06841522, 
    -0.06907488, -0.06794855, -0.06896137, -0.06721681, -0.066843, 
    -0.06709821, -0.06612355, -0.06901795, -0.06789105, -0.07685848, 
    -0.07680228, -0.07654107, -0.0776962, -0.07776748, -0.07884313, 
    -0.07788532, -0.07748107, -0.07646483, -0.07587013, -0.07530928, 
    -0.07409124, -0.07275495, -0.07092833, -0.06964558, -0.06879922, 
    -0.06931695, -0.06885965, -0.06937104, -0.06961212, -0.06698278, 
    -0.06844617, -0.06626283, -0.06638175, -0.0673625, -0.06636833, 
    -0.07676285, -0.07708667, -0.07822181, -0.077332, -0.07896121, 
    -0.07804485, -0.0775229, -0.07554296, -0.07511516, -0.07472054, 
    -0.07394759, -0.0729677, -0.07128113, -0.0698467, -0.06856351, 
    -0.06865671, -0.06862388, -0.06834027, -0.06904495, -0.0682253, 
    -0.06808869, -0.06844641, -0.06639769, -0.06697641, -0.06638428, 
    -0.06676042, -0.07698127, -0.076438, -0.07673106, -0.07618091, 
    -0.07656802, -0.07486203, -0.07435826, -0.07204748, -0.07298683, 
    -0.07149792, -0.07283417, -0.07259548, -0.07144965, -0.07276134, 
    -0.0699249, -0.07183488, -0.06832927, -0.07019109, -0.06821431, 
    -0.06856901, -0.06798284, -0.06746221, -0.06681323, -0.0656326, 
    -0.06590407, -0.06492931, -0.07563553, -0.07494435, -0.07500505, 
    -0.07428822, -0.07376263, -0.07263678, -0.07086805, -0.0715279, 
    -0.07032149, -0.07008183, -0.07191665, -0.07078417, -0.07448553, 
    -0.07387406, -0.07423758, -0.0755807, -0.07137513, -0.07350216, 
    -0.06962456, -0.07073966, -0.06753618, -0.06910992, -0.06605398, 
    -0.06479055, -0.06362492, -0.06228983, -0.07457002, -0.0750365, 
    -0.07420348, -0.07306654, -0.07202812, -0.07067109, -0.07053381, 
    -0.07028303, -0.06963786, -0.06910013, -0.07020383, -0.06896602, 
    -0.07373277, -0.0711936, -0.07521355, -0.0739787, -0.0731331, 
    -0.07350291, -0.07160375, -0.07116356, -0.06940351, -0.07030769, 
    -0.06509994, -0.06735264, -0.0612932, -0.06292703, -0.07520017, 
    -0.07457168, -0.07242629, -0.07343898, -0.07058151, -0.06989598, 
    -0.06934388, -0.06864456, -0.06856958, -0.06815917, -0.06883302, 
    -0.0681857, -0.07066823, -0.06954744, -0.07266837, -0.07189553, 
    -0.07225004, -0.0726409, -0.07144158, -0.07018628, -0.07015988, 
    -0.06976236, -0.06865444, -0.07057017, -0.06481466, -0.06830847, 
    -0.07389253, -0.07270829, -0.07254098, -0.07299623, -0.06996439, 
    -0.07104751, -0.06816917, -0.06893495, -0.0676849, -0.06830309, 
    -0.06839453, -0.06919828, -0.06970359, -0.07099743, -0.07206861, 
    -0.07293005, -0.07272881, -0.07178582, -0.07011028, -0.06856271, 
    -0.06889863, -0.06777907, -0.07078476, -0.0695078, -0.06999843, 
    -0.06872664, -0.07154548, -0.06913716, -0.07217488, -0.07190312, 
    -0.07106919, -0.06942195, -0.06906316, -0.06868188, -0.06891692, 
    -0.07006831, -0.07025892, -0.07108938, -0.07132037, -0.07196221, 
    -0.07249804, -0.07200826, -0.07149757, -0.0700679, -0.06880485, 
    -0.06745481, -0.0671287, -0.0655935, -0.06684019, -0.0647957, 
    -0.06652933, -0.06355829, -0.06900047, -0.06658137, -0.07103154, 
    -0.07053763, -0.06965316, -0.0676682, -0.06873257, -0.06748958, 
    -0.07026642, -0.07175343, -0.07214368, -0.07287733, -0.072127, 
    -0.07218774, -0.07147662, -0.07170435, -0.07002094, -0.07092004, 
    -0.06839678, -0.06749935, -0.06503069, -0.06356389, -0.0621064, 
    -0.06147398, -0.06128285, -0.06120312,
  -0.08618347, -0.08427344, -0.08464142, -0.08312535, -0.08396298, 
    -0.08297516, -0.08579281, -0.08419843, -0.0852128, -0.08600986, 
    -0.08026095, -0.08305837, -0.0774569, -0.07916689, -0.07494235, 
    -0.07772041, -0.07439454, -0.07502125, -0.07315145, -0.07368224, 
    -0.07134189, -0.07290778, -0.07015882, -0.07171282, -0.07146736, 
    -0.07296, -0.08248776, -0.08060391, -0.08260073, -0.08232902, 
    -0.08245087, -0.08394553, -0.08470899, -0.08633139, -0.08603456, 
    -0.08484415, -0.08220714, -0.08309298, -0.08087911, -0.08092845, 
    -0.07853236, -0.07960367, -0.07568386, -0.07677766, -0.07366001, 
    -0.07443175, -0.07369605, -0.07391837, -0.07369316, -0.07482832, 
    -0.07433979, -0.07534669, -0.07940187, -0.07818758, -0.08186588, 
    -0.08416121, -0.08572221, -0.08684752, -0.08668753, -0.08638331, 
    -0.08483724, -0.08340934, -0.08233748, -0.08162826, -0.08093555, 
    -0.07887431, -0.07780537, -0.07546453, -0.07588179, -0.07517641, 
    -0.07450897, -0.07340168, -0.07358281, -0.07309903, -0.07519505, 
    -0.07379529, -0.07612047, -0.07547721, -0.0807476, -0.08285309, 
    -0.08376419, -0.08457053, -0.0865647, -0.08518251, -0.08572468, 
    -0.08444066, -0.08363482, -0.08403243, -0.08160896, -0.08254259, 
    -0.07774247, -0.07977438, -0.07458651, -0.07579597, -0.07429956, 
    -0.07505939, -0.07376219, -0.07492863, -0.07291985, -0.07248967, 
    -0.07278335, -0.07166196, -0.07499382, -0.07369599, -0.08404357, 
    -0.08397858, -0.08367655, -0.08501244, -0.08509489, -0.0863395, 
    -0.08523121, -0.08476359, -0.08358841, -0.08290094, -0.08225279, 
    -0.0808457, -0.07930292, -0.07719567, -0.07571696, -0.07474184, 
    -0.0753383, -0.07481146, -0.07540062, -0.07567841, -0.07265051, 
    -0.07433522, -0.07182217, -0.07195897, -0.07308754, -0.07194354, 
    -0.08393298, -0.08430745, -0.08562052, -0.08459117, -0.08647616, 
    -0.08541577, -0.08481197, -0.08252282, -0.08202848, -0.08157256, 
    -0.0806798, -0.07954848, -0.07760251, -0.07594875, -0.07447036, 
    -0.07457769, -0.07453988, -0.07421325, -0.07502491, -0.07408086, 
    -0.07392354, -0.07433549, -0.0719773, -0.07264318, -0.07196187, 
    -0.07239465, -0.08418556, -0.0835574, -0.08389623, -0.08326018, 
    -0.08370771, -0.08173603, -0.08115409, -0.07848654, -0.07957056, 
    -0.07785257, -0.07939436, -0.07911889, -0.0777969, -0.07931029, 
    -0.07603887, -0.07824127, -0.07420059, -0.0763457, -0.0740682, 
    -0.07447669, -0.07380167, -0.07320231, -0.07245541, -0.07109731, 
    -0.07140951, -0.07028873, -0.08262981, -0.08183113, -0.08190126, 
    -0.08107319, -0.08046622, -0.07916654, -0.07712615, -0.07788714, 
    -0.07649601, -0.07621974, -0.0783356, -0.07702943, -0.08130109, 
    -0.08059489, -0.0810147, -0.08256644, -0.07771094, -0.08016548, 
    -0.07569274, -0.0769781, -0.07328745, -0.07509977, -0.07158194, 
    -0.07012925, -0.06878988, -0.06725694, -0.08139869, -0.0819376, 
    -0.08097532, -0.07966258, -0.0784642, -0.07689905, -0.07674078, 
    -0.07645167, -0.07570808, -0.07508849, -0.07636037, -0.07493399, 
    -0.08043175, -0.07750157, -0.08214217, -0.08071573, -0.07973941, 
    -0.08016634, -0.07797462, -0.07746693, -0.07543802, -0.0764801, 
    -0.07048488, -0.07307618, -0.06611338, -0.06798842, -0.08212671, 
    -0.0814006, -0.07892363, -0.08009252, -0.07679576, -0.07600553, 
    -0.07536931, -0.0745637, -0.07447734, -0.07400471, -0.07478078, 
    -0.07403526, -0.07689575, -0.07560387, -0.07920299, -0.07831123, 
    -0.07872024, -0.07917129, -0.07778757, -0.07634015, -0.07630972, 
    -0.07585155, -0.0745751, -0.0767827, -0.07015696, -0.07417665, 
    -0.08061621, -0.07924908, -0.07905598, -0.07958141, -0.07608438, 
    -0.07733309, -0.07401622, -0.07489821, -0.07345866, -0.07417043, 
    -0.07427573, -0.07520156, -0.07578382, -0.07727535, -0.07851092, 
    -0.07950501, -0.07927274, -0.07818467, -0.07625255, -0.07446943, 
    -0.07485636, -0.07356707, -0.07703011, -0.07555819, -0.07612362, 
    -0.07465825, -0.07790742, -0.07513117, -0.07863352, -0.07831998, 
    -0.07735809, -0.07545927, -0.07504588, -0.07460669, -0.07487743, 
    -0.07620417, -0.07642388, -0.07738137, -0.07764778, -0.07838815, 
    -0.07900643, -0.07844128, -0.07785216, -0.07620369, -0.07474834, 
    -0.07319379, -0.07281844, -0.07105237, -0.07248644, -0.07013517, 
    -0.07212877, -0.06871337, -0.07497368, -0.07218864, -0.07731467, 
    -0.07674518, -0.07572571, -0.07343943, -0.07466508, -0.07323381, 
    -0.07643252, -0.0781473, -0.07859753, -0.07944418, -0.07857829, 
    -0.07864836, -0.077828, -0.07809068, -0.07614957, -0.0771861, 
    -0.07427833, -0.07324505, -0.07040527, -0.0687198, -0.0670464, 
    -0.06632076, -0.0661015, -0.06601005,
  -0.06731972, -0.06577227, -0.0660704, -0.06484208, -0.06552074, 
    -0.06472041, -0.06700322, -0.0657115, -0.06653332, -0.06717906, 
    -0.06252129, -0.06478783, -0.06024928, -0.06163482, -0.05821183, 
    -0.0604628, -0.05776796, -0.05827576, -0.05676073, -0.05719081, 
    -0.05529455, -0.0565633, -0.05433598, -0.05559508, -0.0553962, 
    -0.0566056, -0.06432551, -0.06279916, -0.06441703, -0.06419689, 
    -0.06429562, -0.0655066, -0.06612515, -0.06743955, -0.06719907, 
    -0.06623465, -0.06409815, -0.06481586, -0.06302214, -0.06306211, 
    -0.06112069, -0.06198872, -0.05881265, -0.05969891, -0.0571728, 
    -0.0577981, -0.057202, -0.05738214, -0.05719965, -0.05811943, -0.0577236, 
    -0.05853945, -0.06182522, -0.06084133, -0.06382164, -0.06568135, 
    -0.06694602, -0.06785768, -0.06772807, -0.06748162, -0.06622905, 
    -0.06507218, -0.06420375, -0.06362912, -0.06306786, -0.06139776, 
    -0.06053163, -0.05863493, -0.05897302, -0.05840148, -0.05786068, 
    -0.05696348, -0.05711024, -0.05671826, -0.05841658, -0.05728241, 
    -0.05916642, -0.0586452, -0.06291559, -0.0646215, -0.06535968, 
    -0.06601297, -0.06762857, -0.06650878, -0.06694802, -0.06590775, 
    -0.06525487, -0.065577, -0.06361348, -0.06436993, -0.06048067, 
    -0.06212704, -0.0579235, -0.05890349, -0.057691, -0.05830666, 
    -0.05725559, -0.05820071, -0.05657308, -0.05622452, -0.05646248, 
    -0.05555387, -0.05825353, -0.05720195, -0.06558603, -0.06553337, 
    -0.06528867, -0.06637099, -0.0664378, -0.06744613, -0.06654824, 
    -0.06616938, -0.06521726, -0.06466027, -0.06413513, -0.06299506, 
    -0.06174504, -0.06003761, -0.05883947, -0.05804936, -0.05853265, 
    -0.05810577, -0.05858315, -0.05880823, -0.05635485, -0.05771989, 
    -0.05568368, -0.05579451, -0.05670895, -0.05578202, -0.06549643, 
    -0.06579982, -0.06686363, -0.06602969, -0.06755684, -0.06669775, 
    -0.06620858, -0.06435391, -0.06395338, -0.06358399, -0.06286065, 
    -0.061944, -0.06036727, -0.05902728, -0.05782939, -0.05791636, 
    -0.05788572, -0.05762107, -0.05827872, -0.0575138, -0.05738633, 
    -0.05772011, -0.05580937, -0.0563489, -0.05579687, -0.05614752, 
    -0.06570107, -0.06519213, -0.06546665, -0.06495133, -0.06531392, 
    -0.06371644, -0.06324494, -0.06108356, -0.06196189, -0.06056988, 
    -0.06181912, -0.06159592, -0.06052477, -0.06175101, -0.05910031, 
    -0.06088483, -0.0576108, -0.05934892, -0.05750354, -0.05783452, 
    -0.05728757, -0.05680194, -0.05619676, -0.05509637, -0.05534932, 
    -0.05444123, -0.06444059, -0.0637935, -0.06385031, -0.06317939, 
    -0.06268759, -0.06163453, -0.05998129, -0.06059789, -0.05947071, 
    -0.05924686, -0.06096125, -0.05990292, -0.06336404, -0.06279185, 
    -0.063132, -0.06438926, -0.06045512, -0.06244392, -0.05881985, 
    -0.05986133, -0.05687092, -0.05833938, -0.05548903, -0.05431202, 
    -0.05322686, -0.05198491, -0.06344312, -0.06387975, -0.06310008, 
    -0.06203645, -0.06106545, -0.05979728, -0.05966903, -0.05943478, 
    -0.05883227, -0.05833024, -0.05936081, -0.05820506, -0.06265967, 
    -0.06028548, -0.0640455, -0.06288976, -0.0620987, -0.06244462, 
    -0.06066877, -0.06025741, -0.05861346, -0.05945782, -0.05460016, 
    -0.05669975, -0.05105847, -0.05257753, -0.06403297, -0.06344466, 
    -0.06143771, -0.06238481, -0.05971359, -0.05907329, -0.05855778, 
    -0.05790503, -0.05783504, -0.05745209, -0.05808091, -0.05747684, 
    -0.0597946, -0.05874784, -0.06166407, -0.06094151, -0.06127292, 
    -0.06163838, -0.06051721, -0.05934442, -0.05931976, -0.05894852, 
    -0.05791427, -0.059703, -0.05433448, -0.05759142, -0.06280912, 
    -0.06170142, -0.06154495, -0.06197068, -0.05913718, -0.06014897, 
    -0.05746142, -0.05817606, -0.05700964, -0.05758637, -0.05767169, 
    -0.05842186, -0.05889364, -0.06010218, -0.06110331, -0.06190878, 
    -0.06172058, -0.06083897, -0.05927344, -0.05782864, -0.05814215, 
    -0.05709749, -0.05990347, -0.05871083, -0.05916897, -0.05798163, 
    -0.06061432, -0.05836483, -0.06120265, -0.0609486, -0.06016922, 
    -0.05863068, -0.05829572, -0.05793986, -0.05815922, -0.05923424, 
    -0.05941226, -0.06018808, -0.06040395, -0.06100384, -0.0615048, 
    -0.06104689, -0.06056955, -0.05923385, -0.05805463, -0.05679503, 
    -0.05649091, -0.05505996, -0.05622191, -0.05431682, -0.05593212, 
    -0.05316487, -0.05823722, -0.05598062, -0.06013404, -0.05967261, 
    -0.05884656, -0.05699407, -0.05798716, -0.05682747, -0.05941926, 
    -0.06080869, -0.06117349, -0.06185949, -0.06115789, -0.06121467, 
    -0.06054997, -0.06076281, -0.05919, -0.06002986, -0.0576738, -0.05683657, 
    -0.05453566, -0.05317007, -0.05181434, -0.05122647, -0.05104884, 
    -0.05097475,
  -0.06391447, -0.06222166, -0.06254755, -0.06120564, -0.06194681, 
    -0.06107282, -0.06356799, -0.06215525, -0.0630538, -0.06376047, 
    -0.05867587, -0.06114641, -0.05620678, -0.0577116, -0.0539992, 
    -0.05643849, -0.05351913, -0.05406837, -0.05243093, -0.05289538, 
    -0.05084988, -0.05221782, -0.04981819, -0.05117367, -0.05095939, 
    -0.05226349, -0.0606419, -0.05897837, -0.06074176, -0.0605016, 
    -0.06060929, -0.06193136, -0.06260741, -0.06404568, -0.06378238, 
    -0.06272715, -0.0603939, -0.06117702, -0.05922118, -0.05926472, 
    -0.05715287, -0.05809643, -0.05464952, -0.05560982, -0.05287593, 
    -0.05355172, -0.05290747, -0.0531021, -0.05290494, -0.05389924, 
    -0.05347117, -0.05435374, -0.05791861, -0.05684945, -0.06009239, 
    -0.0621223, -0.06350538, -0.0645037, -0.0643617, -0.06409176, 
    -0.06272102, -0.06145686, -0.06050907, -0.05988252, -0.05927098, 
    -0.05745393, -0.05651321, -0.0544571, -0.0548232, -0.05420442, 
    -0.05361939, -0.05264986, -0.05280836, -0.05238508, -0.05422076, 
    -0.05299434, -0.0550327, -0.05446822, -0.05910514, -0.06096487, 
    -0.06177086, -0.06248477, -0.0642527, -0.06302696, -0.06350757, 
    -0.06236975, -0.06165637, -0.06200828, -0.05986547, -0.06069036, 
    -0.05645789, -0.05824688, -0.05368733, -0.05474789, -0.05343593, 
    -0.05410181, -0.05296537, -0.05398717, -0.05222838, -0.0518523, 
    -0.05210903, -0.05112926, -0.05404432, -0.05290742, -0.06201814, 
    -0.06196061, -0.06169329, -0.06287625, -0.06294931, -0.06405289, 
    -0.06307013, -0.06265578, -0.0616153, -0.06100719, -0.06043423, 
    -0.05919169, -0.05783143, -0.05597714, -0.05467856, -0.05382345, 
    -0.05434638, -0.05388446, -0.05440104, -0.05464473, -0.05199289, 
    -0.05346716, -0.05126915, -0.05138862, -0.05237504, -0.05137514, 
    -0.06192025, -0.06225177, -0.06341521, -0.06250305, -0.06417414, 
    -0.0632337, -0.06269864, -0.06067289, -0.06023603, -0.05983333, 
    -0.05904532, -0.05804779, -0.05633481, -0.05488196, -0.05358555, 
    -0.0536796, -0.05364647, -0.05336033, -0.05407158, -0.05324438, 
    -0.05310663, -0.0534674, -0.05140464, -0.05198648, -0.05139116, 
    -0.05176925, -0.06214385, -0.06158786, -0.06188772, -0.06132491, 
    -0.06172087, -0.0599777, -0.05946387, -0.05711254, -0.05806725, 
    -0.05655472, -0.05791198, -0.05766932, -0.05650576, -0.05783793, 
    -0.05496107, -0.05689669, -0.05334923, -0.05523045, -0.0532333, 
    -0.05359109, -0.05299992, -0.05247543, -0.05182235, -0.05063646, 
    -0.05090889, -0.04993139, -0.06076746, -0.0600617, -0.06012364, 
    -0.05939246, -0.0588569, -0.05771129, -0.05591604, -0.05658513, 
    -0.05536243, -0.05511985, -0.05697969, -0.05583104, -0.05959363, 
    -0.05897041, -0.05934083, -0.06071145, -0.05643016, -0.05859167, 
    -0.05465731, -0.05578594, -0.05254991, -0.05413722, -0.0510594, 
    -0.04979242, -0.04862646, -0.04729465, -0.0596798, -0.06015574, 
    -0.05930608, -0.05814834, -0.05709287, -0.05571648, -0.05557742, 
    -0.05532349, -0.05467076, -0.05412732, -0.05524332, -0.05399187, 
    -0.05882651, -0.05624605, -0.06033648, -0.05907702, -0.05821606, 
    -0.05859243, -0.05666208, -0.05621559, -0.05443385, -0.05534846, 
    -0.05010237, -0.05236511, -0.04630303, -0.0479298, -0.06032282, 
    -0.05968148, -0.05749736, -0.05852734, -0.05562573, -0.05493181, 
    -0.05437358, -0.05366734, -0.05359167, -0.0531777, -0.05385758, 
    -0.05320444, -0.05571358, -0.05457934, -0.0577434, -0.05695825, 
    -0.05731827, -0.05771548, -0.05649755, -0.05522557, -0.05519884, 
    -0.05479667, -0.05367734, -0.05561425, -0.04981658, -0.05332828, 
    -0.05898922, -0.05778401, -0.05761391, -0.05807681, -0.05500102, 
    -0.05609793, -0.05318778, -0.0539605, -0.05269971, -0.05332283, 
    -0.05341506, -0.05422647, -0.05473723, -0.05604718, -0.05713399, 
    -0.05800948, -0.05780485, -0.05684688, -0.05514865, -0.05358474, 
    -0.05392382, -0.05279458, -0.05583163, -0.05453927, -0.05503546, 
    -0.05375019, -0.05660297, -0.05416476, -0.05724192, -0.05696594, 
    -0.05611991, -0.05445249, -0.05408997, -0.05370501, -0.05394229, 
    -0.05510618, -0.05529909, -0.05614037, -0.05637461, -0.05702594, 
    -0.05757027, -0.05707271, -0.05655436, -0.05510575, -0.05382914, 
    -0.05246797, -0.05213971, -0.05059725, -0.05184948, -0.04979759, 
    -0.05153696, -0.04855993, -0.05402667, -0.05158925, -0.05608174, 
    -0.0555813, -0.05468624, -0.05268289, -0.05375617, -0.05250299, 
    -0.05530667, -0.056814, -0.05721024, -0.05795588, -0.05719329, 
    -0.05725498, -0.0565331, -0.05676418, -0.05505824, -0.05596872, 
    -0.05341733, -0.05251282, -0.05003298, -0.04856551, -0.04711195, 
    -0.04648273, -0.04629274, -0.04621351,
  -0.04035198, -0.03907359, -0.03931955, -0.03830725, -0.03886621, 
    -0.03820712, -0.04009016, -0.03902347, -0.03970177, -0.0402356, 
    -0.03640241, -0.03826259, -0.03454811, -0.03567765, -0.03289467, 
    -0.03472191, -0.0325357, -0.03294641, -0.03172283, -0.03206963, 
    -0.03054395, -0.03156378, -0.02977613, -0.03078516, -0.03062552, 
    -0.03159786, -0.03788236, -0.03662992, -0.0379576, -0.03777665, 
    -0.03785779, -0.03885455, -0.03936473, -0.04045115, -0.04025215, 
    -0.03945512, -0.03769551, -0.03828567, -0.0368126, -0.03684536, 
    -0.03525804, -0.0359668, -0.03338129, -0.03410057, -0.03205509, 
    -0.03256006, -0.03207865, -0.03222404, -0.03207676, -0.03281991, 
    -0.03249985, -0.03315991, -0.03583318, -0.03503027, -0.03746841, 
    -0.03899861, -0.04004287, -0.0407974, -0.04069003, -0.04048597, 
    -0.0394505, -0.03849666, -0.03778228, -0.03731038, -0.03685007, 
    -0.03548411, -0.03477797, -0.03323727, -0.03351131, -0.03304819, 
    -0.03261065, -0.03188627, -0.03200463, -0.03168861, -0.03306041, 
    -0.03214354, -0.03366819, -0.03324559, -0.03672529, -0.03812575, 
    -0.03873348, -0.03927216, -0.04060763, -0.0396815, -0.04004452, 
    -0.03918534, -0.03864712, -0.03891259, -0.03729754, -0.03791887, 
    -0.03473647, -0.03607988, -0.03266144, -0.03345493, -0.0324735, 
    -0.03297142, -0.0321219, -0.03288567, -0.03157166, -0.03129108, 
    -0.0314826, -0.03075207, -0.03292842, -0.03207862, -0.03892003, 
    -0.03887662, -0.03867497, -0.0395677, -0.03962287, -0.04045659, 
    -0.0397141, -0.03940124, -0.03861614, -0.03815764, -0.03772589, 
    -0.03679041, -0.03576767, -0.03437591, -0.03340303, -0.03276323, 
    -0.03315441, -0.03280886, -0.03319531, -0.03337771, -0.03139596, 
    -0.03249685, -0.03085631, -0.03094536, -0.03168111, -0.03093531, 
    -0.03884617, -0.03909631, -0.03997475, -0.03928595, -0.04054824, 
    -0.03983764, -0.0394336, -0.03790571, -0.0375766, -0.03727334, 
    -0.03668029, -0.03593025, -0.03464414, -0.03355532, -0.03258535, 
    -0.03265566, -0.03263089, -0.032417, -0.03294881, -0.03233036, 
    -0.03222743, -0.03249703, -0.03095729, -0.03139117, -0.03094725, 
    -0.03122914, -0.03901487, -0.03859545, -0.03882163, -0.03839717, 
    -0.03869577, -0.03738204, -0.03699523, -0.03522776, -0.03594487, 
    -0.03480911, -0.0358282, -0.03564588, -0.03477238, -0.03577255, 
    -0.03361456, -0.03506573, -0.03240871, -0.03381631, -0.03232207, 
    -0.0325895, -0.03214771, -0.03175604, -0.03126875, -0.03038502, 
    -0.0305879, -0.02986032, -0.03797697, -0.0374453, -0.03749195, 
    -0.03694149, -0.03653856, -0.03567741, -0.03433011, -0.03483192, 
    -0.03391519, -0.03373347, -0.03512803, -0.03426639, -0.0370929, 
    -0.03662394, -0.03690264, -0.03793476, -0.03471566, -0.03633909, 
    -0.03338712, -0.03423258, -0.03181165, -0.03299791, -0.03070002, 
    -0.02975696, -0.02889069, -0.02790317, -0.03715776, -0.03751612, 
    -0.03687648, -0.03600582, -0.03521299, -0.03418051, -0.03407629, 
    -0.03388602, -0.03339719, -0.03299051, -0.03382596, -0.03288919, 
    -0.0365157, -0.03457757, -0.03765226, -0.03670414, -0.03605671, 
    -0.03633966, -0.03488967, -0.03455472, -0.03321987, -0.03390472, 
    -0.02998751, -0.0316737, -0.02716934, -0.02837385, -0.03764197, 
    -0.03715903, -0.03551672, -0.03629072, -0.03411249, -0.03359264, 
    -0.03317476, -0.0326465, -0.03258992, -0.03228053, -0.03278875, 
    -0.03230051, -0.03417834, -0.03332876, -0.03570153, -0.03511194, 
    -0.03538223, -0.03568055, -0.03476622, -0.03381266, -0.03379264, 
    -0.03349145, -0.03265397, -0.03410389, -0.02977493, -0.03239306, 
    -0.03663808, -0.03573204, -0.03560426, -0.03595205, -0.03364447, 
    -0.03446649, -0.03228806, -0.03286572, -0.03192349, -0.03238898, 
    -0.03245791, -0.03306468, -0.03344695, -0.03442843, -0.03524387, 
    -0.03590146, -0.0357477, -0.03502835, -0.03375505, -0.03258475, 
    -0.03283829, -0.03199434, -0.03426683, -0.03329876, -0.03367027, 
    -0.03270845, -0.03484531, -0.03301851, -0.0353249, -0.03511771, 
    -0.03448297, -0.03323382, -0.03296256, -0.03267466, -0.0328521, 
    -0.03372323, -0.03386774, -0.03449832, -0.034674, -0.03516275, 
    -0.03557148, -0.03519786, -0.03480884, -0.03372291, -0.03276749, 
    -0.03175048, -0.03150549, -0.03035583, -0.03128898, -0.02976081, 
    -0.03105594, -0.02884131, -0.03291522, -0.03109493, -0.03445435, 
    -0.03407919, -0.03340878, -0.03191093, -0.03271292, -0.03177662, 
    -0.03387342, -0.03500367, -0.03530111, -0.03586118, -0.03528839, 
    -0.0353347, -0.03479289, -0.03496628, -0.03368732, -0.03436961, 
    -0.03245961, -0.03178396, -0.02993588, -0.02884545, -0.02776788, 
    -0.02730223, -0.02716173, -0.02710316,
  -0.01970498, -0.01870054, -0.01889315, -0.01810236, -0.01853836, 
    -0.01802443, -0.01949861, -0.01866132, -0.0191931, -0.01961321, 
    -0.01662923, -0.0180676, -0.01521544, -0.01607415, -0.01397336, 
    -0.01534705, -0.01370618, -0.01401194, -0.01310463, -0.01336067, 
    -0.01224115, -0.0129875, -0.01168477, -0.01241693, -0.01230054, 
    -0.01301258, -0.01777204, -0.01680411, -0.01783047, -0.01769001, 
    -0.01775297, -0.01852925, -0.01892857, -0.01978323, -0.01962626, 
    -0.01899946, -0.01762709, -0.01808556, -0.01694474, -0.01696998, 
    -0.01575423, -0.01629523, -0.01433699, -0.01487744, -0.01334993, 
    -0.01372429, -0.01336735, -0.01347497, -0.01336595, -0.01391764, 
    -0.01367955, -0.01417136, -0.016193, -0.01558102, -0.01745117, 
    -0.01864188, -0.01946137, -0.02005681, -0.01997192, -0.01981072, 
    -0.01899583, -0.01824993, -0.01769438, -0.01732891, -0.01697361, 
    -0.01592645, -0.01538954, -0.0142292, -0.01443443, -0.0140879, 
    -0.01376189, -0.01322518, -0.01331261, -0.01307941, -0.01409703, 
    -0.01341536, -0.01455215, -0.01423542, -0.01687751, -0.01796114, 
    -0.01843468, -0.01885602, -0.0199068, -0.01917717, -0.01946267, 
    -0.01878802, -0.01836728, -0.01857461, -0.01731899, -0.01780039, 
    -0.01535808, -0.01638183, -0.01379967, -0.01439216, -0.01365998, 
    -0.0140306, -0.01339934, -0.01396665, -0.0129933, -0.01278713, 
    -0.01292779, -0.01239279, -0.01399853, -0.01336732, -0.01858043, 
    -0.0185465, -0.01838901, -0.0190878, -0.01913112, -0.01978753, 
    -0.01920278, -0.0189572, -0.01834311, -0.01798595, -0.01765065, 
    -0.01692765, -0.01614293, -0.01508524, -0.01435328, -0.01387542, 
    -0.01416725, -0.0139094, -0.01419783, -0.01433431, -0.01286412, 
    -0.01367732, -0.01246887, -0.01253393, -0.01307388, -0.01252659, 
    -0.01852271, -0.01871832, -0.01940775, -0.01886683, -0.01985989, 
    -0.01929989, -0.01898258, -0.01779017, -0.01753494, -0.01730028, 
    -0.01684286, -0.01626726, -0.01528814, -0.01446743, -0.01374308, 
    -0.01379537, -0.01377694, -0.01361804, -0.01401373, -0.01355376, 
    -0.01347748, -0.01367746, -0.01254266, -0.0128606, -0.01253532, 
    -0.0127417, -0.01865459, -0.01832696, -0.01850353, -0.01817239, 
    -0.01840525, -0.01738434, -0.01708553, -0.01573118, -0.01627845, 
    -0.01541315, -0.0161892, -0.01604989, -0.0153853, -0.01614666, 
    -0.01451188, -0.01560796, -0.01361189, -0.01466344, -0.01354762, 
    -0.01374616, -0.01341845, -0.01312911, -0.01277074, -0.01212558, 
    -0.01227314, -0.01174553, -0.01784551, -0.01743328, -0.01746939, 
    -0.01704408, -0.01673384, -0.01607397, -0.01505064, -0.01543046, 
    -0.01473782, -0.01460118, -0.01565532, -0.01500252, -0.0171609, 
    -0.01679951, -0.01701413, -0.01781273, -0.01534232, -0.01658061, 
    -0.01434136, -0.014977, -0.01317011, -0.01405037, -0.01235483, 
    -0.01167095, -0.01104943, -0.01034922, -0.01721098, -0.0174881, 
    -0.01699397, -0.0163251, -0.01571995, -0.01493772, -0.01485914, 
    -0.01471587, -0.0143489, -0.01404485, -0.0146707, -0.01396927, 
    -0.01671627, -0.01523773, -0.01759356, -0.01686122, -0.01636408, 
    -0.01658105, -0.01547426, -0.01522044, -0.01421619, -0.01472995, 
    -0.01183745, -0.01306842, -0.009834968, -0.01068182, -0.01758559, 
    -0.01721196, -0.01595132, -0.01654349, -0.01488643, -0.01449544, 
    -0.01418246, -0.01378855, -0.01374648, -0.01351682, -0.01389443, 
    -0.01353163, -0.01493608, -0.01429766, -0.0160924, -0.01564309, 
    -0.0158488, -0.01607637, -0.01538063, -0.0146607, -0.01464565, 
    -0.01441954, -0.01379411, -0.01487995, -0.0116839, -0.01360027, 
    -0.01681039, -0.0161157, -0.01601812, -0.01628395, -0.01453434, 
    -0.0151537, -0.0135224, -0.01395178, -0.01325267, -0.01359724, 
    -0.0136484, -0.01410022, -0.01438618, -0.01512493, -0.01574344, 
    -0.01624523, -0.01612766, -0.01557956, -0.01461739, -0.01374263, 
    -0.01393133, -0.01330501, -0.01500286, -0.01427521, -0.01455371, 
    -0.01383464, -0.01544061, -0.01406575, -0.01580513, -0.01564748, 
    -0.01516616, -0.01422662, -0.014024, -0.0138095, -0.01394163, 
    -0.01459348, -0.01470212, -0.01517777, -0.01531075, -0.01568172, 
    -0.0159931, -0.01570843, -0.01541295, -0.01459324, -0.01387859, 
    -0.01312501, -0.01294462, -0.01210438, -0.01278559, -0.01167372, 
    -0.01261482, -0.01101419, -0.01398868, -0.01264336, -0.01514452, 
    -0.01486133, -0.01435758, -0.0132434, -0.01383797, -0.01314428, 
    -0.01470639, -0.01556082, -0.01578701, -0.01621442, -0.01577733, 
    -0.0158126, -0.01540086, -0.01553242, -0.01456652, -0.01508047, 
    -0.01364966, -0.01314969, -0.01180012, -0.01101715, -0.01025401, 
    -0.009927695, -0.009829662, -0.009788851,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15 ;

 SOILWATER_10CM =
  297.8986, 299.1539, 298.9096, 299.9243, 299.3612, 300.0261, 298.1528, 
    299.2037, 298.5326, 298.0115, 301.9005, 299.9697, 303.8941, 302.6757, 
    305.7423, 303.7043, 306.1546, 305.6836, 307.1034, 306.6961, 308.5174, 
    307.2915, 309.4651, 308.2244, 308.4182, 307.2511, 300.3578, 301.6601, 
    300.2808, 300.4662, 300.383, 299.3727, 298.8645, 297.8029, 297.9955, 
    298.7753, 300.5496, 299.9465, 301.4686, 301.4341, 303.1251, 302.3652, 
    305.1902, 304.3869, 306.7131, 306.1268, 306.6855, 306.5161, 306.6877, 
    305.8282, 306.1962, 305.4407, 302.5084, 303.3703, 300.7841, 299.2282, 
    298.1988, 297.4699, 297.5728, 297.7692, 298.7799, 299.7328, 300.4606, 
    300.9482, 301.4292, 302.8824, 303.6435, 305.3528, 305.0439, 305.5674, 
    306.0685, 306.9109, 306.7721, 307.1437, 305.5538, 306.6096, 304.8681, 
    305.3436, 301.5594, 300.1091, 299.4938, 298.9565, 297.652, 298.5523, 
    298.1971, 299.0428, 299.5811, 299.3148, 300.9615, 300.3205, 303.6887, 
    302.2441, 306.01, 305.1073, 306.2267, 305.6552, 306.6349, 305.7531, 
    307.2821, 307.6158, 307.3877, 308.2647, 305.7042, 306.6855, 299.3073, 
    299.3508, 299.5532, 298.6643, 298.61, 297.7976, 298.5205, 298.8286, 
    299.6124, 300.0766, 300.5185, 301.4918, 302.5786, 304.083, 305.1658, 
    305.8932, 305.4471, 305.8409, 305.4006, 305.1945, 307.4907, 306.1996, 
    308.1385, 308.0309, 307.1525, 308.0431, 299.3813, 299.1315, 298.2653, 
    298.943, 297.7093, 298.3993, 298.7965, 300.3337, 300.6724, 300.9866, 
    301.6079, 302.4043, 303.7895, 304.9944, 306.0977, 306.0168, 306.0452, 
    306.292, 305.6809, 306.3925, 306.5119, 306.1995, 308.0165, 307.4966, 
    308.0287, 307.69, 299.2127, 299.6332, 299.4059, 299.8334, 299.5321, 
    300.8734, 301.2765, 303.1573, 302.3886, 303.6098, 302.5138, 302.71, 
    303.6492, 302.5737, 304.9277, 303.3317, 306.3016, 304.7019, 306.4021, 
    306.0929, 306.605, 307.0641, 307.6426, 308.7121, 308.4642, 309.3604, 
    300.261, 300.808, 300.7599, 301.3332, 301.7574, 302.6761, 304.1335, 
    303.5853, 304.5925, 304.795, 303.2651, 304.2036, 301.1746, 301.6671, 
    301.3739, 300.3041, 303.7114, 301.9682, 305.1837, 304.241, 306.9986, 
    305.6246, 308.3278, 309.4887, 310.585, 311.8693, 301.107, 300.7349, 
    301.4015, 302.3232, 303.1735, 304.2984, 304.4138, 304.6249, 305.1725, 
    305.6334, 304.6916, 305.749, 301.7808, 303.8621, 300.5942, 301.5824, 
    302.2689, 301.9679, 303.5227, 303.8874, 305.3726, 304.6042, 309.2018, 
    307.161, 312.8504, 311.2522, 300.605, 301.1057, 302.8481, 302.0198, 
    304.3737, 304.9526, 305.424, 306.0271, 306.0924, 306.4503, 305.864, 
    306.4271, 304.3008, 305.2496, 302.6502, 303.2823, 302.9921, 302.6728, 
    303.6567, 304.7063, 304.729, 305.0661, 306.0173, 304.3832, 309.4655, 
    306.3187, 301.6525, 302.6169, 302.755, 302.381, 304.8945, 303.9839, 
    306.4416, 305.7758, 306.8672, 306.3245, 306.2447, 305.549, 305.1163, 
    304.0255, 303.1403, 302.4353, 302.6005, 303.3724, 304.7707, 306.0982, 
    305.807, 306.7842, 304.2033, 305.2834, 304.8655, 305.956, 303.5707, 
    305.6003, 303.0535, 303.2762, 303.9658, 305.3566, 305.6653, 305.9947, 
    305.7914, 304.8063, 304.6452, 303.9491, 303.757, 303.2277, 302.79, 
    303.1898, 303.6102, 304.8068, 305.8882, 307.0706, 307.3607, 308.7473, 
    307.6178, 309.4831, 307.8963, 310.6474, 305.7186, 307.8501, 303.9973, 
    304.4106, 305.159, 306.8815, 305.9509, 307.0396, 304.6389, 303.3989, 
    303.079, 302.4784, 303.0927, 303.043, 303.6277, 303.4398, 304.8466, 
    304.0903, 306.2427, 307.031, 309.2663, 310.6426, 312.0489, 312.6712, 
    312.8608, 312.9401 ;

 SOMC_FIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOMHR =
  6.357484e-08, 6.385439e-08, 6.380004e-08, 6.402553e-08, 6.390044e-08, 
    6.404809e-08, 6.363151e-08, 6.386549e-08, 6.371612e-08, 6.360001e-08, 
    6.446311e-08, 6.403558e-08, 6.490716e-08, 6.463451e-08, 6.53194e-08, 
    6.486474e-08, 6.541108e-08, 6.530627e-08, 6.562168e-08, 6.553132e-08, 
    6.593476e-08, 6.566339e-08, 6.614388e-08, 6.586995e-08, 6.59128e-08, 
    6.565443e-08, 6.412161e-08, 6.440989e-08, 6.410454e-08, 6.414565e-08, 
    6.41272e-08, 6.390303e-08, 6.379007e-08, 6.355347e-08, 6.359642e-08, 
    6.377019e-08, 6.416413e-08, 6.40304e-08, 6.436741e-08, 6.43598e-08, 
    6.473498e-08, 6.456582e-08, 6.519642e-08, 6.501719e-08, 6.55351e-08, 
    6.540485e-08, 6.552898e-08, 6.549134e-08, 6.552947e-08, 6.533845e-08, 
    6.542029e-08, 6.52522e-08, 6.459751e-08, 6.478992e-08, 6.421605e-08, 
    6.387099e-08, 6.364178e-08, 6.347913e-08, 6.350213e-08, 6.354596e-08, 
    6.377121e-08, 6.398299e-08, 6.414438e-08, 6.425233e-08, 6.43587e-08, 
    6.46807e-08, 6.48511e-08, 6.523266e-08, 6.51638e-08, 6.528045e-08, 
    6.539189e-08, 6.557899e-08, 6.55482e-08, 6.563063e-08, 6.527737e-08, 
    6.551215e-08, 6.512457e-08, 6.523057e-08, 6.438765e-08, 6.406648e-08, 
    6.392999e-08, 6.38105e-08, 6.351981e-08, 6.372055e-08, 6.364142e-08, 
    6.382967e-08, 6.39493e-08, 6.389013e-08, 6.425529e-08, 6.411333e-08, 
    6.48612e-08, 6.453907e-08, 6.537889e-08, 6.517793e-08, 6.542706e-08, 
    6.529993e-08, 6.551776e-08, 6.532171e-08, 6.566131e-08, 6.573526e-08, 
    6.568472e-08, 6.587883e-08, 6.531085e-08, 6.552898e-08, 6.388848e-08, 
    6.389813e-08, 6.394308e-08, 6.374548e-08, 6.373339e-08, 6.355229e-08, 
    6.371343e-08, 6.378205e-08, 6.395624e-08, 6.405927e-08, 6.415721e-08, 
    6.437256e-08, 6.461306e-08, 6.494936e-08, 6.519095e-08, 6.53529e-08, 
    6.525359e-08, 6.534127e-08, 6.524326e-08, 6.519733e-08, 6.570755e-08, 
    6.542106e-08, 6.585091e-08, 6.582712e-08, 6.563259e-08, 6.582981e-08, 
    6.390491e-08, 6.384938e-08, 6.365659e-08, 6.380746e-08, 6.353257e-08, 
    6.368644e-08, 6.377493e-08, 6.41163e-08, 6.41913e-08, 6.426085e-08, 
    6.43982e-08, 6.457448e-08, 6.488371e-08, 6.515276e-08, 6.539837e-08, 
    6.538038e-08, 6.538671e-08, 6.544158e-08, 6.530567e-08, 6.546389e-08, 
    6.549045e-08, 6.542102e-08, 6.582394e-08, 6.570883e-08, 6.582662e-08, 
    6.575167e-08, 6.386743e-08, 6.396086e-08, 6.391037e-08, 6.400531e-08, 
    6.393843e-08, 6.423585e-08, 6.432501e-08, 6.474225e-08, 6.457101e-08, 
    6.484353e-08, 6.459869e-08, 6.464208e-08, 6.485244e-08, 6.461192e-08, 
    6.513793e-08, 6.478133e-08, 6.544371e-08, 6.508762e-08, 6.546603e-08, 
    6.539731e-08, 6.551109e-08, 6.561299e-08, 6.574118e-08, 6.597772e-08, 
    6.592295e-08, 6.612076e-08, 6.410015e-08, 6.422135e-08, 6.421067e-08, 
    6.433749e-08, 6.443128e-08, 6.463457e-08, 6.496062e-08, 6.483801e-08, 
    6.506309e-08, 6.510828e-08, 6.476632e-08, 6.497628e-08, 6.430245e-08, 
    6.441132e-08, 6.434649e-08, 6.410971e-08, 6.486627e-08, 6.447801e-08, 
    6.519495e-08, 6.498462e-08, 6.559846e-08, 6.529319e-08, 6.589279e-08, 
    6.614913e-08, 6.639036e-08, 6.667229e-08, 6.428748e-08, 6.420513e-08, 
    6.435257e-08, 6.455657e-08, 6.474583e-08, 6.499745e-08, 6.502319e-08, 
    6.507033e-08, 6.519242e-08, 6.529509e-08, 6.508524e-08, 6.532083e-08, 
    6.443658e-08, 6.489997e-08, 6.4174e-08, 6.439262e-08, 6.454454e-08, 
    6.44779e-08, 6.482399e-08, 6.490557e-08, 6.523705e-08, 6.506569e-08, 
    6.608587e-08, 6.563452e-08, 6.688694e-08, 6.653695e-08, 6.417636e-08, 
    6.428719e-08, 6.467292e-08, 6.448939e-08, 6.501424e-08, 6.514343e-08, 
    6.524845e-08, 6.538271e-08, 6.53972e-08, 6.547674e-08, 6.53464e-08, 
    6.547159e-08, 6.499798e-08, 6.520963e-08, 6.462883e-08, 6.47702e-08, 
    6.470516e-08, 6.463382e-08, 6.485399e-08, 6.508855e-08, 6.509355e-08, 
    6.516876e-08, 6.538072e-08, 6.501637e-08, 6.614414e-08, 6.544767e-08, 
    6.440805e-08, 6.462153e-08, 6.465201e-08, 6.456932e-08, 6.513049e-08, 
    6.492716e-08, 6.54748e-08, 6.532679e-08, 6.55693e-08, 6.544879e-08, 
    6.543107e-08, 6.527629e-08, 6.517993e-08, 6.493648e-08, 6.473839e-08, 
    6.458131e-08, 6.461784e-08, 6.479039e-08, 6.51029e-08, 6.539852e-08, 
    6.533376e-08, 6.555087e-08, 6.497619e-08, 6.521717e-08, 6.512403e-08, 
    6.536688e-08, 6.483475e-08, 6.528791e-08, 6.471893e-08, 6.476881e-08, 
    6.492312e-08, 6.523352e-08, 6.530218e-08, 6.537551e-08, 6.533025e-08, 
    6.511083e-08, 6.507487e-08, 6.491937e-08, 6.487644e-08, 6.475795e-08, 
    6.465985e-08, 6.474948e-08, 6.48436e-08, 6.511091e-08, 6.535181e-08, 
    6.561444e-08, 6.567871e-08, 6.598559e-08, 6.573579e-08, 6.614802e-08, 
    6.579756e-08, 6.640422e-08, 6.531416e-08, 6.578724e-08, 6.493014e-08, 
    6.502248e-08, 6.518949e-08, 6.557254e-08, 6.536574e-08, 6.560759e-08, 
    6.507346e-08, 6.479635e-08, 6.472464e-08, 6.459086e-08, 6.472769e-08, 
    6.471657e-08, 6.48475e-08, 6.480542e-08, 6.511979e-08, 6.495092e-08, 
    6.543063e-08, 6.560568e-08, 6.610003e-08, 6.640308e-08, 6.671156e-08, 
    6.684775e-08, 6.68892e-08, 6.690653e-08 ;

 SOM_C_LEACHED =
  4.487101e-20, 4.254831e-20, -1.960332e-20, 1.69865e-20, 4.408414e-20, 
    -2.441936e-21, 4.624704e-20, 2.53491e-21, -1.984593e-20, -3.18578e-20, 
    -1.532834e-20, 3.814324e-20, -1.933366e-20, -3.104988e-20, -2.775303e-20, 
    8.909278e-22, -3.637645e-20, 6.506488e-20, -6.140348e-20, 4.540946e-21, 
    9.452574e-21, 1.770222e-20, 2.189577e-20, -6.424227e-20, 1.752194e-20, 
    -4.13449e-21, -5.062767e-20, -1.163998e-22, 5.883461e-20, 1.554555e-20, 
    6.558239e-21, 8.575249e-21, -1.348952e-20, 5.486501e-21, 2.348061e-20, 
    4.148553e-20, 2.908582e-22, -5.686385e-21, -4.959846e-20, -1.587094e-21, 
    -1.354382e-21, -5.537999e-21, -1.0647e-20, 4.543079e-20, 4.667087e-20, 
    -1.60037e-21, 5.961247e-21, 2.745358e-20, 5.370867e-21, 3.646423e-21, 
    1.767861e-21, 1.906789e-20, 5.89056e-20, -1.632877e-20, 1.269569e-20, 
    2.948089e-20, -2.059322e-20, -6.221669e-20, -2.914325e-20, 1.999523e-20, 
    -4.426142e-20, 1.983043e-20, -2.68553e-20, -4.823551e-20, -2.647139e-20, 
    -9.221046e-21, -3.343311e-20, 2.549176e-20, 4.892866e-20, 6.870198e-21, 
    3.835959e-20, 1.811119e-20, 2.400238e-20, 3.129297e-21, -7.462809e-21, 
    6.034398e-20, 7.647472e-20, 4.164882e-21, 2.994305e-20, 2.509464e-20, 
    3.605328e-20, -2.166756e-20, -3.333096e-20, 6.443891e-20, -1.940709e-20, 
    -9.341227e-21, 3.29385e-20, -1.799918e-21, 4.238617e-20, -3.830725e-20, 
    -3.953297e-21, 3.556853e-20, -1.575771e-20, -1.877288e-20, 4.723183e-21, 
    -1.592931e-21, -7.473624e-20, -1.404487e-21, 3.066776e-20, -5.043399e-20, 
    4.939473e-20, -4.039831e-20, -1.95051e-20, 5.41797e-21, -3.36739e-20, 
    -5.507423e-20, 6.907831e-21, -1.140863e-20, 5.495071e-20, 5.577674e-21, 
    -4.162326e-21, -5.758657e-21, 2.908099e-20, 2.119914e-20, -2.122647e-20, 
    -1.687452e-20, -3.779948e-20, -2.251708e-20, 3.420466e-20, 2.138746e-20, 
    -9.027614e-21, 7.763581e-20, -2.175812e-21, 1.049276e-19, -4.548571e-20, 
    5.11663e-20, 1.63712e-20, 5.353148e-20, 9.137922e-20, -1.178408e-20, 
    9.379658e-21, 2.723912e-20, -3.463669e-21, 2.170861e-20, -3.274884e-20, 
    2.221454e-20, -1.870936e-20, -5.760157e-20, 6.257405e-20, 4.774296e-20, 
    4.632131e-20, 2.195783e-20, -1.226704e-20, 5.539177e-21, 7.154248e-21, 
    -8.342735e-20, -4.750856e-20, 1.974566e-20, -1.772318e-20, -9.425545e-21, 
    7.185643e-21, 8.588153e-21, 4.702569e-21, -7.654394e-20, 3.335577e-20, 
    2.069734e-20, -3.490141e-20, 3.682177e-20, 1.485224e-20, -5.204346e-20, 
    -4.516797e-20, 8.411146e-21, 7.161389e-22, 5.246985e-20, 4.943066e-20, 
    3.454084e-20, -1.815557e-20, -3.218347e-20, 3.27738e-20, -2.840668e-20, 
    3.243152e-21, -7.705389e-21, 1.085245e-20, 3.957974e-20, -2.658849e-20, 
    1.181348e-20, 4.886824e-20, 3.531267e-21, 6.087366e-20, -2.840815e-20, 
    -7.803239e-20, 2.426984e-20, 5.457809e-21, -4.585277e-20, -7.410932e-21, 
    1.083215e-20, 3.666794e-20, -2.26547e-20, 1.895428e-20, -2.850359e-21, 
    7.903097e-20, -1.856021e-20, 8.910258e-20, -5.497237e-20, -5.194889e-20, 
    -2.220937e-20, 1.745732e-20, 7.223696e-21, 5.793782e-20, -1.391063e-20, 
    1.75233e-20, -1.218823e-20, -8.281423e-21, 3.547674e-20, 3.239202e-20, 
    -2.99842e-20, 6.545352e-20, 6.147654e-20, -8.234326e-20, 1.325186e-21, 
    -2.3307e-20, -2.547414e-20, 5.079844e-20, -9.340347e-21, -8.319893e-21, 
    -9.547479e-21, -3.103584e-21, 3.568432e-20, 4.333487e-20, 1.746441e-20, 
    -4.916035e-20, 8.369034e-22, -5.449302e-21, 1.701911e-20, 1.932823e-20, 
    3.860409e-20, 1.250401e-21, -9.728994e-20, -5.705605e-20, -2.584818e-21, 
    1.609842e-20, -3.181067e-20, 2.444346e-20, -7.888318e-21, 6.300314e-21, 
    9.042932e-21, -7.875753e-20, -2.054242e-20, -7.074812e-20, -2.728585e-20, 
    6.868994e-21, -1.353735e-20, 4.83821e-20, -4.060544e-20, -5.939053e-21, 
    -6.048461e-22, -6.745268e-20, 2.232163e-20, -5.298515e-20, 8.125703e-21, 
    2.478611e-20, 3.237949e-20, -6.562965e-20, 9.087546e-21, -3.25307e-20, 
    4.977072e-20, -2.704297e-20, 1.880039e-20, 2.808033e-21, -2.763486e-20, 
    3.705918e-20, -1.58539e-20, -1.033383e-19, 2.300674e-21, -4.57082e-20, 
    2.852323e-20, -8.358281e-20, -5.157016e-21, -6.744847e-20, -9.663643e-21, 
    4.05518e-20, -1.341966e-20, 1.311714e-20, 2.55261e-21, 6.807174e-20, 
    -2.974418e-20, -6.326483e-20, -4.977429e-22, -1.403602e-20, 
    -5.157159e-21, -1.472741e-20, -1.149146e-20, 2.285982e-20, 2.795566e-21, 
    -2.131886e-20, 1.900533e-21, 4.583892e-21, -1.525229e-20, 7.735222e-20, 
    -1.336115e-20, 6.334725e-20, 5.023534e-20, 5.783399e-20, -3.207679e-20, 
    3.530376e-20, -5.576083e-20, -1.33946e-20, -9.91963e-21, -2.794462e-20, 
    -3.875302e-20, 4.566681e-21, -2.296542e-20, -2.711215e-20, -1.686223e-22, 
    7.258363e-20, 1.403177e-20, 4.853781e-20, -2.155094e-20, -3.245391e-20, 
    3.759104e-20, -9.999427e-22, 2.838115e-20, -2.354333e-20, 4.545935e-20, 
    -1.379925e-20, -2.873991e-20, 7.187448e-21, 1.053225e-20, 3.516349e-20, 
    4.062966e-20, -4.555978e-20, -4.988311e-20, -2.632616e-20, 1.855082e-20, 
    1.114179e-20, 9.04854e-21, 2.040469e-20, -9.077144e-20, 1.096886e-20, 
    8.558356e-20, 4.019558e-20, -5.575147e-20, 2.307911e-20, -5.690389e-20, 
    -3.61156e-20, 1.053613e-19, -7.653055e-21, 2.608118e-20 ;

 SR =
  6.35757e-08, 6.385525e-08, 6.38009e-08, 6.402639e-08, 6.39013e-08, 
    6.404895e-08, 6.363237e-08, 6.386636e-08, 6.371699e-08, 6.360087e-08, 
    6.446398e-08, 6.403645e-08, 6.490803e-08, 6.463537e-08, 6.532027e-08, 
    6.48656e-08, 6.541195e-08, 6.530715e-08, 6.562256e-08, 6.55322e-08, 
    6.593564e-08, 6.566426e-08, 6.614476e-08, 6.587083e-08, 6.591368e-08, 
    6.565531e-08, 6.412248e-08, 6.441076e-08, 6.41054e-08, 6.41465e-08, 
    6.412806e-08, 6.390389e-08, 6.379094e-08, 6.355432e-08, 6.359728e-08, 
    6.377105e-08, 6.416499e-08, 6.403126e-08, 6.436827e-08, 6.436066e-08, 
    6.473585e-08, 6.456669e-08, 6.519728e-08, 6.501806e-08, 6.553597e-08, 
    6.540572e-08, 6.552985e-08, 6.549221e-08, 6.553034e-08, 6.533932e-08, 
    6.542116e-08, 6.525307e-08, 6.459837e-08, 6.479079e-08, 6.421691e-08, 
    6.387185e-08, 6.364264e-08, 6.347999e-08, 6.350298e-08, 6.354682e-08, 
    6.377208e-08, 6.398385e-08, 6.414524e-08, 6.42532e-08, 6.435957e-08, 
    6.468156e-08, 6.485197e-08, 6.523354e-08, 6.516466e-08, 6.528133e-08, 
    6.539276e-08, 6.557987e-08, 6.554907e-08, 6.563151e-08, 6.527824e-08, 
    6.551303e-08, 6.512544e-08, 6.523145e-08, 6.438852e-08, 6.406734e-08, 
    6.393085e-08, 6.381136e-08, 6.352067e-08, 6.372141e-08, 6.364228e-08, 
    6.383054e-08, 6.395017e-08, 6.3891e-08, 6.425615e-08, 6.411419e-08, 
    6.486207e-08, 6.453993e-08, 6.537977e-08, 6.51788e-08, 6.542793e-08, 
    6.53008e-08, 6.551863e-08, 6.532259e-08, 6.566219e-08, 6.573613e-08, 
    6.56856e-08, 6.587971e-08, 6.531172e-08, 6.552985e-08, 6.388935e-08, 
    6.389899e-08, 6.394394e-08, 6.374634e-08, 6.373425e-08, 6.355315e-08, 
    6.371429e-08, 6.378291e-08, 6.39571e-08, 6.406013e-08, 6.415808e-08, 
    6.437342e-08, 6.461393e-08, 6.495023e-08, 6.519183e-08, 6.535377e-08, 
    6.525447e-08, 6.534214e-08, 6.524414e-08, 6.519819e-08, 6.570843e-08, 
    6.542193e-08, 6.585179e-08, 6.5828e-08, 6.563347e-08, 6.583068e-08, 
    6.390577e-08, 6.385024e-08, 6.365745e-08, 6.380832e-08, 6.353343e-08, 
    6.36873e-08, 6.377579e-08, 6.411717e-08, 6.419216e-08, 6.426171e-08, 
    6.439907e-08, 6.457535e-08, 6.488458e-08, 6.515364e-08, 6.539925e-08, 
    6.538125e-08, 6.538759e-08, 6.544246e-08, 6.530654e-08, 6.546477e-08, 
    6.549133e-08, 6.542189e-08, 6.582482e-08, 6.570971e-08, 6.58275e-08, 
    6.575254e-08, 6.386828e-08, 6.396172e-08, 6.391124e-08, 6.400618e-08, 
    6.393929e-08, 6.423671e-08, 6.432588e-08, 6.474312e-08, 6.457188e-08, 
    6.484441e-08, 6.459956e-08, 6.464295e-08, 6.485331e-08, 6.461279e-08, 
    6.513881e-08, 6.47822e-08, 6.544459e-08, 6.508849e-08, 6.546691e-08, 
    6.539818e-08, 6.551196e-08, 6.561386e-08, 6.574206e-08, 6.59786e-08, 
    6.592382e-08, 6.612164e-08, 6.410102e-08, 6.422221e-08, 6.421153e-08, 
    6.433836e-08, 6.443215e-08, 6.463544e-08, 6.496149e-08, 6.483888e-08, 
    6.506396e-08, 6.510916e-08, 6.476719e-08, 6.497716e-08, 6.430331e-08, 
    6.441219e-08, 6.434736e-08, 6.411058e-08, 6.486714e-08, 6.447888e-08, 
    6.519582e-08, 6.498549e-08, 6.559934e-08, 6.529407e-08, 6.589367e-08, 
    6.615002e-08, 6.639124e-08, 6.667317e-08, 6.428834e-08, 6.4206e-08, 
    6.435344e-08, 6.455743e-08, 6.47467e-08, 6.499832e-08, 6.502406e-08, 
    6.507121e-08, 6.51933e-08, 6.529596e-08, 6.508611e-08, 6.53217e-08, 
    6.443745e-08, 6.490084e-08, 6.417487e-08, 6.439348e-08, 6.454541e-08, 
    6.447876e-08, 6.482487e-08, 6.490644e-08, 6.523793e-08, 6.506657e-08, 
    6.608675e-08, 6.56354e-08, 6.688783e-08, 6.653783e-08, 6.417723e-08, 
    6.428806e-08, 6.467379e-08, 6.449026e-08, 6.501512e-08, 6.514431e-08, 
    6.524932e-08, 6.538358e-08, 6.539807e-08, 6.547761e-08, 6.534727e-08, 
    6.547247e-08, 6.499886e-08, 6.52105e-08, 6.46297e-08, 6.477106e-08, 
    6.470603e-08, 6.463469e-08, 6.485485e-08, 6.508942e-08, 6.509442e-08, 
    6.516963e-08, 6.53816e-08, 6.501724e-08, 6.614502e-08, 6.544855e-08, 
    6.440892e-08, 6.462241e-08, 6.465289e-08, 6.457019e-08, 6.513136e-08, 
    6.492802e-08, 6.547567e-08, 6.532767e-08, 6.557018e-08, 6.544967e-08, 
    6.543194e-08, 6.527716e-08, 6.51808e-08, 6.493735e-08, 6.473926e-08, 
    6.458218e-08, 6.46187e-08, 6.479126e-08, 6.510376e-08, 6.539939e-08, 
    6.533463e-08, 6.555175e-08, 6.497706e-08, 6.521804e-08, 6.512491e-08, 
    6.536776e-08, 6.483562e-08, 6.528879e-08, 6.471979e-08, 6.476968e-08, 
    6.492399e-08, 6.52344e-08, 6.530306e-08, 6.537638e-08, 6.533113e-08, 
    6.51117e-08, 6.507574e-08, 6.492024e-08, 6.487731e-08, 6.475882e-08, 
    6.466072e-08, 6.475035e-08, 6.484448e-08, 6.511178e-08, 6.535268e-08, 
    6.561532e-08, 6.567959e-08, 6.598647e-08, 6.573666e-08, 6.61489e-08, 
    6.579844e-08, 6.64051e-08, 6.531504e-08, 6.578811e-08, 6.493101e-08, 
    6.502334e-08, 6.519036e-08, 6.557342e-08, 6.536661e-08, 6.560847e-08, 
    6.507433e-08, 6.479721e-08, 6.47255e-08, 6.459173e-08, 6.472857e-08, 
    6.471743e-08, 6.484837e-08, 6.480629e-08, 6.512066e-08, 6.49518e-08, 
    6.54315e-08, 6.560656e-08, 6.610091e-08, 6.640397e-08, 6.671245e-08, 
    6.684864e-08, 6.689009e-08, 6.690742e-08 ;

 STORVEGC =
  0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545 ;

 STORVEGN =
  0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061 ;

 SUPPLEMENT_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SoilAlpha =
  0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 
    0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999934, 0.9999933, 
    0.9999934, 0.9999934, 0.9999935, 0.9999934, 0.9999935, 0.9999935, 
    0.9999935, 0.9999935, 0.9999936, 0.9999935, 0.9999936, 0.9999936, 
    0.9999936, 0.9999935, 0.9999933, 0.9999934, 0.9999933, 0.9999933, 
    0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 
    0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 
    0.9999935, 0.9999935, 0.9999935, 0.9999934, 0.9999934, 0.9999934, 
    0.9999933, 0.9999933, 0.9999933, 0.9999932, 0.9999932, 0.9999933, 
    0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999935, 0.9999935, 
    0.9999935, 0.9999935, 0.9999934, 0.9999935, 0.9999934, 0.9999934, 
    0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999932, 0.9999933, 
    0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 
    0.9999934, 0.9999934, 0.9999935, 0.9999934, 0.9999935, 0.9999935, 
    0.9999935, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 0.9999936, 
    0.9999935, 0.9999935, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 
    0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 
    0.9999933, 0.9999933, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 
    0.9999934, 0.9999935, 0.9999934, 0.9999934, 0.9999935, 0.9999935, 
    0.9999936, 0.9999936, 0.9999935, 0.9999936, 0.9999933, 0.9999933, 
    0.9999933, 0.9999933, 0.9999932, 0.9999933, 0.9999933, 0.9999933, 
    0.9999933, 0.9999933, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999935, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 
    0.9999935, 0.9999935, 0.9999936, 0.9999935, 0.9999936, 0.9999936, 
    0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 
    0.9999933, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999934, 
    0.9999935, 0.9999935, 0.9999935, 0.9999935, 0.9999936, 0.9999936, 
    0.9999936, 0.9999936, 0.9999933, 0.9999933, 0.9999933, 0.9999933, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999933, 0.9999934, 0.9999933, 0.9999933, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999935, 
    0.9999936, 0.9999936, 0.9999936, 0.9999936, 0.9999933, 0.9999933, 
    0.9999933, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999935, 0.9999934, 0.9999935, 0.9999934, 0.9999934, 
    0.9999933, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999936, 0.9999935, 0.9999937, 0.9999936, 
    0.9999933, 0.9999933, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999934, 
    0.9999936, 0.9999935, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999935, 0.9999935, 0.9999935, 0.9999935, 
    0.9999935, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999935, 0.9999935, 
    0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999934, 0.9999935, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999935, 
    0.9999935, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 0.9999935, 
    0.9999935, 0.9999936, 0.9999935, 0.9999936, 0.9999936, 0.9999936, 
    0.9999935, 0.9999936, 0.9999934, 0.9999934, 0.9999934, 0.9999935, 
    0.9999935, 0.9999935, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 0.9999934, 
    0.9999935, 0.9999935, 0.9999936, 0.9999936, 0.9999937, 0.9999937, 
    0.9999937, 0.9999937 ;

 SoilAlpha_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TAUX =
  -0.1477094, -0.1477245, -0.1477216, -0.1477333, -0.147727, -0.1477344, 
    -0.1477125, -0.147725, -0.1477171, -0.1477109, -0.1477537, -0.1477338, 
    -0.1477685, -0.1477599, -0.1477925, -0.1477671, -0.1477954, -0.1477923, 
    -0.1478021, -0.1477993, -0.1478115, -0.1478034, -0.1478181, -0.1478097, 
    -0.1478109, -0.1478031, -0.1477383, -0.1477517, -0.1477374, -0.1477394, 
    -0.1477386, -0.1477271, -0.1477208, -0.1477084, -0.1477107, -0.1477199, 
    -0.1477403, -0.1477337, -0.1477508, -0.1477504, -0.1477632, -0.1477577, 
    -0.1477889, -0.147772, -0.1477994, -0.1477954, -0.1477992, -0.1477981, 
    -0.1477992, -0.1477933, -0.1477958, -0.1477906, -0.1477587, -0.147765, 
    -0.147743, -0.147725, -0.1477131, -0.1477043, -0.1477056, -0.1477079, 
    -0.1477199, -0.1477313, -0.1477395, -0.1477449, -0.1477503, -0.1477611, 
    -0.1477668, -0.1477899, -0.1477879, -0.1477914, -0.147795, -0.1478007, 
    -0.1477998, -0.1478023, -0.1477914, -0.1477986, -0.1477753, -0.14779, 
    -0.1477509, -0.1477356, -0.1477282, -0.1477221, -0.1477065, -0.1477172, 
    -0.147713, -0.1477233, -0.1477296, -0.1477266, -0.1477451, -0.1477379, 
    -0.1477671, -0.1477567, -0.1477946, -0.1477883, -0.1477961, -0.1477921, 
    -0.1477988, -0.1477928, -0.1478033, -0.1478055, -0.147804, -0.1478101, 
    -0.1477925, -0.1477992, -0.1477264, -0.1477269, -0.1477294, -0.1477186, 
    -0.147718, -0.1477083, -0.147717, -0.1477206, -0.14773, -0.1477352, 
    -0.1477401, -0.1477509, -0.1477591, -0.1477698, -0.1477887, -0.1477938, 
    -0.1477907, -0.1477934, -0.1477904, -0.147789, -0.1478046, -0.1477958, 
    -0.1478092, -0.1478085, -0.1478024, -0.1478085, -0.1477273, -0.1477244, 
    -0.1477139, -0.1477221, -0.1477072, -0.1477154, -0.1477201, -0.1477379, 
    -0.1477419, -0.1477453, -0.1477519, -0.147758, -0.1477679, -0.1477875, 
    -0.1477952, -0.1477946, -0.1477948, -0.1477965, -0.1477923, -0.1477972, 
    -0.147798, -0.1477959, -0.1478084, -0.1478048, -0.1478084, -0.1478061, 
    -0.1477253, -0.1477302, -0.1477276, -0.1477324, -0.147729, -0.1477439, 
    -0.1477483, -0.1477633, -0.1477578, -0.1477666, -0.1477588, -0.1477602, 
    -0.1477667, -0.1477592, -0.1477869, -0.1477645, -0.1477966, -0.1477738, 
    -0.1477973, -0.1477952, -0.1477987, -0.1478018, -0.1478058, -0.147813, 
    -0.1478114, -0.1478175, -0.1477373, -0.1477432, -0.1477429, -0.1477492, 
    -0.147753, -0.14776, -0.1477702, -0.1477666, -0.1477734, -0.1477747, 
    -0.1477643, -0.1477707, -0.1477473, -0.1477521, -0.1477496, -0.1477376, 
    -0.1477673, -0.1477546, -0.1477888, -0.147771, -0.1478013, -0.1477918, 
    -0.1478104, -0.1478181, -0.1478259, -0.1478343, -0.1477467, -0.1477426, 
    -0.14775, -0.1477572, -0.1477636, -0.1477713, -0.1477722, -0.1477736, 
    -0.1477888, -0.147792, -0.1477739, -0.1477928, -0.1477528, -0.1477684, 
    -0.1477409, -0.1477514, -0.1477569, -0.1477547, -0.1477662, -0.1477686, 
    -0.1477901, -0.1477735, -0.1478161, -0.1478023, -0.1478412, -0.1478302, 
    -0.1477411, -0.1477467, -0.1477611, -0.1477552, -0.1477719, -0.1477872, 
    -0.1477906, -0.1477946, -0.1477951, -0.1477976, -0.1477936, -0.1477975, 
    -0.1477714, -0.1477893, -0.1477598, -0.1477644, -0.1477623, -0.14776, 
    -0.1477671, -0.147774, -0.1477743, -0.147788, -0.147794, -0.147772, 
    -0.1478176, -0.1477962, -0.1477522, -0.1477593, -0.1477605, -0.1477579, 
    -0.1477754, -0.1477692, -0.1477975, -0.147793, -0.1478005, -0.1477967, 
    -0.1477962, -0.1477914, -0.1477884, -0.1477695, -0.1477633, -0.1477583, 
    -0.1477595, -0.147765, -0.1477744, -0.1477951, -0.1477931, -0.1477999, 
    -0.1477707, -0.1477895, -0.1477751, -0.1477942, -0.1477665, -0.1477912, 
    -0.1477628, -0.1477644, -0.1477691, -0.1477899, -0.1477922, -0.1477944, 
    -0.1477931, -0.1477747, -0.1477737, -0.147769, -0.1477677, -0.1477641, 
    -0.1477608, -0.1477637, -0.1477667, -0.1477748, -0.1477937, -0.1478018, 
    -0.1478039, -0.147813, -0.1478053, -0.1478177, -0.1478068, -0.1478258, 
    -0.1477922, -0.1478069, -0.1477694, -0.1477722, -0.1477885, -0.1478004, 
    -0.1477942, -0.1478015, -0.1477737, -0.1477651, -0.147763, -0.1477585, 
    -0.147763, -0.1477627, -0.1477669, -0.1477656, -0.1477751, -0.14777, 
    -0.1477961, -0.1478015, -0.1478168, -0.1478261, -0.1478358, -0.14784, 
    -0.1478413, -0.1478418 ;

 TAUY =
  -0.1477094, -0.1477245, -0.1477216, -0.1477333, -0.147727, -0.1477344, 
    -0.1477125, -0.147725, -0.1477171, -0.1477109, -0.1477537, -0.1477338, 
    -0.1477685, -0.1477599, -0.1477925, -0.1477671, -0.1477954, -0.1477923, 
    -0.1478021, -0.1477993, -0.1478115, -0.1478034, -0.1478181, -0.1478097, 
    -0.1478109, -0.1478031, -0.1477383, -0.1477517, -0.1477374, -0.1477394, 
    -0.1477386, -0.1477271, -0.1477208, -0.1477084, -0.1477107, -0.1477199, 
    -0.1477403, -0.1477337, -0.1477508, -0.1477504, -0.1477632, -0.1477577, 
    -0.1477889, -0.147772, -0.1477994, -0.1477954, -0.1477992, -0.1477981, 
    -0.1477992, -0.1477933, -0.1477958, -0.1477906, -0.1477587, -0.147765, 
    -0.147743, -0.147725, -0.1477131, -0.1477043, -0.1477056, -0.1477079, 
    -0.1477199, -0.1477313, -0.1477395, -0.1477449, -0.1477503, -0.1477611, 
    -0.1477668, -0.1477899, -0.1477879, -0.1477914, -0.147795, -0.1478007, 
    -0.1477998, -0.1478023, -0.1477914, -0.1477986, -0.1477753, -0.14779, 
    -0.1477509, -0.1477356, -0.1477282, -0.1477221, -0.1477065, -0.1477172, 
    -0.147713, -0.1477233, -0.1477296, -0.1477266, -0.1477451, -0.1477379, 
    -0.1477671, -0.1477567, -0.1477946, -0.1477883, -0.1477961, -0.1477921, 
    -0.1477988, -0.1477928, -0.1478033, -0.1478055, -0.147804, -0.1478101, 
    -0.1477925, -0.1477992, -0.1477264, -0.1477269, -0.1477294, -0.1477186, 
    -0.147718, -0.1477083, -0.147717, -0.1477206, -0.14773, -0.1477352, 
    -0.1477401, -0.1477509, -0.1477591, -0.1477698, -0.1477887, -0.1477938, 
    -0.1477907, -0.1477934, -0.1477904, -0.147789, -0.1478046, -0.1477958, 
    -0.1478092, -0.1478085, -0.1478024, -0.1478085, -0.1477273, -0.1477244, 
    -0.1477139, -0.1477221, -0.1477072, -0.1477154, -0.1477201, -0.1477379, 
    -0.1477419, -0.1477453, -0.1477519, -0.147758, -0.1477679, -0.1477875, 
    -0.1477952, -0.1477946, -0.1477948, -0.1477965, -0.1477923, -0.1477972, 
    -0.147798, -0.1477959, -0.1478084, -0.1478048, -0.1478084, -0.1478061, 
    -0.1477253, -0.1477302, -0.1477276, -0.1477324, -0.147729, -0.1477439, 
    -0.1477483, -0.1477633, -0.1477578, -0.1477666, -0.1477588, -0.1477602, 
    -0.1477667, -0.1477592, -0.1477869, -0.1477645, -0.1477966, -0.1477738, 
    -0.1477973, -0.1477952, -0.1477987, -0.1478018, -0.1478058, -0.147813, 
    -0.1478114, -0.1478175, -0.1477373, -0.1477432, -0.1477429, -0.1477492, 
    -0.147753, -0.14776, -0.1477702, -0.1477666, -0.1477734, -0.1477747, 
    -0.1477643, -0.1477707, -0.1477473, -0.1477521, -0.1477496, -0.1477376, 
    -0.1477673, -0.1477546, -0.1477888, -0.147771, -0.1478013, -0.1477918, 
    -0.1478104, -0.1478181, -0.1478259, -0.1478343, -0.1477467, -0.1477426, 
    -0.14775, -0.1477572, -0.1477636, -0.1477713, -0.1477722, -0.1477736, 
    -0.1477888, -0.147792, -0.1477739, -0.1477928, -0.1477528, -0.1477684, 
    -0.1477409, -0.1477514, -0.1477569, -0.1477547, -0.1477662, -0.1477686, 
    -0.1477901, -0.1477735, -0.1478161, -0.1478023, -0.1478412, -0.1478302, 
    -0.1477411, -0.1477467, -0.1477611, -0.1477552, -0.1477719, -0.1477872, 
    -0.1477906, -0.1477946, -0.1477951, -0.1477976, -0.1477936, -0.1477975, 
    -0.1477714, -0.1477893, -0.1477598, -0.1477644, -0.1477623, -0.14776, 
    -0.1477671, -0.147774, -0.1477743, -0.147788, -0.147794, -0.147772, 
    -0.1478176, -0.1477962, -0.1477522, -0.1477593, -0.1477605, -0.1477579, 
    -0.1477754, -0.1477692, -0.1477975, -0.147793, -0.1478005, -0.1477967, 
    -0.1477962, -0.1477914, -0.1477884, -0.1477695, -0.1477633, -0.1477583, 
    -0.1477595, -0.147765, -0.1477744, -0.1477951, -0.1477931, -0.1477999, 
    -0.1477707, -0.1477895, -0.1477751, -0.1477942, -0.1477665, -0.1477912, 
    -0.1477628, -0.1477644, -0.1477691, -0.1477899, -0.1477922, -0.1477944, 
    -0.1477931, -0.1477747, -0.1477737, -0.147769, -0.1477677, -0.1477641, 
    -0.1477608, -0.1477637, -0.1477667, -0.1477748, -0.1477937, -0.1478018, 
    -0.1478039, -0.147813, -0.1478053, -0.1478177, -0.1478068, -0.1478258, 
    -0.1477922, -0.1478069, -0.1477694, -0.1477722, -0.1477885, -0.1478004, 
    -0.1477942, -0.1478015, -0.1477737, -0.1477651, -0.147763, -0.1477585, 
    -0.147763, -0.1477627, -0.1477669, -0.1477656, -0.1477751, -0.14777, 
    -0.1477961, -0.1478015, -0.1478168, -0.1478261, -0.1478358, -0.14784, 
    -0.1478413, -0.1478418 ;

 TBOT =
  256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044 ;

 TBUILD =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TG =
  262.7732, 262.7871, 262.7844, 262.7957, 262.7894, 262.7968, 262.7761, 
    262.7877, 262.7803, 262.7745, 262.8174, 262.7961, 262.8397, 262.8261, 
    262.8603, 262.8376, 262.8649, 262.8596, 262.8755, 262.8709, 262.8911, 
    262.8776, 262.9016, 262.8879, 262.89, 262.8771, 262.8004, 262.8148, 
    262.7996, 262.8016, 262.8007, 262.7896, 262.7839, 262.7722, 262.7743, 
    262.7829, 262.8026, 262.7959, 262.8127, 262.8123, 262.8311, 262.8226, 
    262.8541, 262.8453, 262.8711, 262.8646, 262.8708, 262.8689, 262.8708, 
    262.8612, 262.8654, 262.8569, 262.8242, 262.8339, 262.8051, 262.7879, 
    262.7766, 262.7685, 262.7696, 262.7718, 262.783, 262.7935, 262.8016, 
    262.807, 262.8123, 262.8283, 262.8369, 262.8559, 262.8525, 262.8583, 
    262.8639, 262.8733, 262.8718, 262.8759, 262.8582, 262.87, 262.8506, 
    262.8558, 262.8136, 262.7977, 262.7909, 262.7849, 262.7705, 262.7805, 
    262.7766, 262.7859, 262.7919, 262.7889, 262.8071, 262.8, 262.8374, 
    262.8213, 262.8633, 262.8532, 262.8657, 262.8593, 262.8702, 262.8604, 
    262.8774, 262.8811, 262.8786, 262.8884, 262.8599, 262.8708, 262.7888, 
    262.7893, 262.7916, 262.7817, 262.7811, 262.7721, 262.7801, 262.7835, 
    262.7922, 262.7973, 262.8022, 262.813, 262.825, 262.8419, 262.8539, 
    262.862, 262.857, 262.8614, 262.8565, 262.8542, 262.8798, 262.8654, 
    262.887, 262.8858, 262.876, 262.8859, 262.7896, 262.7869, 262.7773, 
    262.7848, 262.7711, 262.7788, 262.7832, 262.8002, 262.8039, 262.8074, 
    262.8142, 262.8231, 262.8386, 262.8519, 262.8643, 262.8633, 262.8637, 
    262.8664, 262.8596, 262.8676, 262.8689, 262.8654, 262.8856, 262.8798, 
    262.8857, 262.882, 262.7878, 262.7924, 262.7899, 262.7946, 262.7913, 
    262.8061, 262.8105, 262.8315, 262.8229, 262.8365, 262.8243, 262.8264, 
    262.8369, 262.825, 262.8512, 262.8334, 262.8665, 262.8488, 262.8676, 
    262.8642, 262.8699, 262.875, 262.8814, 262.8933, 262.8906, 262.9005, 
    262.7994, 262.8054, 262.8049, 262.8112, 262.8159, 262.8261, 262.8424, 
    262.8363, 262.8476, 262.8498, 262.8327, 262.8432, 262.8094, 262.8149, 
    262.8116, 262.7998, 262.8377, 262.8182, 262.854, 262.8436, 262.8743, 
    262.8589, 262.8891, 262.9019, 262.914, 262.9281, 262.8087, 262.8046, 
    262.812, 262.8221, 262.8316, 262.8443, 262.8456, 262.8479, 262.8539, 
    262.8591, 262.8487, 262.8604, 262.8161, 262.8394, 262.803, 262.8139, 
    262.8216, 262.8182, 262.8356, 262.8397, 262.8561, 262.8477, 262.8987, 
    262.8761, 262.9389, 262.9214, 262.8032, 262.8087, 262.828, 262.8188, 
    262.8451, 262.8515, 262.8567, 262.8635, 262.8642, 262.8682, 262.8616, 
    262.8679, 262.8443, 262.8548, 262.8258, 262.8329, 262.8296, 262.826, 
    262.8371, 262.8488, 262.8491, 262.8527, 262.8633, 262.8452, 262.9016, 
    262.8666, 262.8147, 262.8254, 262.8269, 262.8228, 262.851, 262.8407, 
    262.8681, 262.8607, 262.8728, 262.8668, 262.8659, 262.8581, 262.8533, 
    262.8412, 262.8313, 262.8234, 262.8253, 262.8339, 262.8495, 262.8643, 
    262.861, 262.8719, 262.8432, 262.8552, 262.8506, 262.8627, 262.8361, 
    262.8586, 262.8303, 262.8328, 262.8405, 262.856, 262.8594, 262.8631, 
    262.8608, 262.8499, 262.8481, 262.8404, 262.8382, 262.8323, 262.8274, 
    262.8318, 262.8365, 262.85, 262.8619, 262.8751, 262.8783, 262.8937, 
    262.8811, 262.9018, 262.8842, 262.9147, 262.86, 262.8837, 262.8409, 
    262.8455, 262.8538, 262.873, 262.8626, 262.8747, 262.8481, 262.8342, 
    262.8306, 262.8239, 262.8307, 262.8302, 262.8368, 262.8347, 262.8504, 
    262.8419, 262.8659, 262.8746, 262.8994, 262.9146, 262.9301, 262.937, 
    262.9391, 262.9399 ;

 TG_R =
  262.7732, 262.7871, 262.7844, 262.7957, 262.7894, 262.7968, 262.7761, 
    262.7877, 262.7803, 262.7745, 262.8174, 262.7961, 262.8397, 262.8261, 
    262.8603, 262.8376, 262.8649, 262.8596, 262.8755, 262.8709, 262.8911, 
    262.8776, 262.9016, 262.8879, 262.89, 262.8771, 262.8004, 262.8148, 
    262.7996, 262.8016, 262.8007, 262.7896, 262.7839, 262.7722, 262.7743, 
    262.7829, 262.8026, 262.7959, 262.8127, 262.8123, 262.8311, 262.8226, 
    262.8541, 262.8453, 262.8711, 262.8646, 262.8708, 262.8689, 262.8708, 
    262.8612, 262.8654, 262.8569, 262.8242, 262.8339, 262.8051, 262.7879, 
    262.7766, 262.7685, 262.7696, 262.7718, 262.783, 262.7935, 262.8016, 
    262.807, 262.8123, 262.8283, 262.8369, 262.8559, 262.8525, 262.8583, 
    262.8639, 262.8733, 262.8718, 262.8759, 262.8582, 262.87, 262.8506, 
    262.8558, 262.8136, 262.7977, 262.7909, 262.7849, 262.7705, 262.7805, 
    262.7766, 262.7859, 262.7919, 262.7889, 262.8071, 262.8, 262.8374, 
    262.8213, 262.8633, 262.8532, 262.8657, 262.8593, 262.8702, 262.8604, 
    262.8774, 262.8811, 262.8786, 262.8884, 262.8599, 262.8708, 262.7888, 
    262.7893, 262.7916, 262.7817, 262.7811, 262.7721, 262.7801, 262.7835, 
    262.7922, 262.7973, 262.8022, 262.813, 262.825, 262.8419, 262.8539, 
    262.862, 262.857, 262.8614, 262.8565, 262.8542, 262.8798, 262.8654, 
    262.887, 262.8858, 262.876, 262.8859, 262.7896, 262.7869, 262.7773, 
    262.7848, 262.7711, 262.7788, 262.7832, 262.8002, 262.8039, 262.8074, 
    262.8142, 262.8231, 262.8386, 262.8519, 262.8643, 262.8633, 262.8637, 
    262.8664, 262.8596, 262.8676, 262.8689, 262.8654, 262.8856, 262.8798, 
    262.8857, 262.882, 262.7878, 262.7924, 262.7899, 262.7946, 262.7913, 
    262.8061, 262.8105, 262.8315, 262.8229, 262.8365, 262.8243, 262.8264, 
    262.8369, 262.825, 262.8512, 262.8334, 262.8665, 262.8488, 262.8676, 
    262.8642, 262.8699, 262.875, 262.8814, 262.8933, 262.8906, 262.9005, 
    262.7994, 262.8054, 262.8049, 262.8112, 262.8159, 262.8261, 262.8424, 
    262.8363, 262.8476, 262.8498, 262.8327, 262.8432, 262.8094, 262.8149, 
    262.8116, 262.7998, 262.8377, 262.8182, 262.854, 262.8436, 262.8743, 
    262.8589, 262.8891, 262.9019, 262.914, 262.9281, 262.8087, 262.8046, 
    262.812, 262.8221, 262.8316, 262.8443, 262.8456, 262.8479, 262.8539, 
    262.8591, 262.8487, 262.8604, 262.8161, 262.8394, 262.803, 262.8139, 
    262.8216, 262.8182, 262.8356, 262.8397, 262.8561, 262.8477, 262.8987, 
    262.8761, 262.9389, 262.9214, 262.8032, 262.8087, 262.828, 262.8188, 
    262.8451, 262.8515, 262.8567, 262.8635, 262.8642, 262.8682, 262.8616, 
    262.8679, 262.8443, 262.8548, 262.8258, 262.8329, 262.8296, 262.826, 
    262.8371, 262.8488, 262.8491, 262.8527, 262.8633, 262.8452, 262.9016, 
    262.8666, 262.8147, 262.8254, 262.8269, 262.8228, 262.851, 262.8407, 
    262.8681, 262.8607, 262.8728, 262.8668, 262.8659, 262.8581, 262.8533, 
    262.8412, 262.8313, 262.8234, 262.8253, 262.8339, 262.8495, 262.8643, 
    262.861, 262.8719, 262.8432, 262.8552, 262.8506, 262.8627, 262.8361, 
    262.8586, 262.8303, 262.8328, 262.8405, 262.856, 262.8594, 262.8631, 
    262.8608, 262.8499, 262.8481, 262.8404, 262.8382, 262.8323, 262.8274, 
    262.8318, 262.8365, 262.85, 262.8619, 262.8751, 262.8783, 262.8937, 
    262.8811, 262.9018, 262.8842, 262.9147, 262.86, 262.8837, 262.8409, 
    262.8455, 262.8538, 262.873, 262.8626, 262.8747, 262.8481, 262.8342, 
    262.8306, 262.8239, 262.8307, 262.8302, 262.8368, 262.8347, 262.8504, 
    262.8419, 262.8659, 262.8746, 262.8994, 262.9146, 262.9301, 262.937, 
    262.9391, 262.9399 ;

 TG_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TH2OSFC =
  255.0004, 255, 255.0001, 254.9997, 254.9999, 254.9997, 255.0003, 255, 
    255.0002, 255.0004, 254.9991, 254.9997, 254.9985, 254.9989, 254.9979, 
    254.9985, 254.9978, 254.998, 254.9976, 254.9977, 254.9972, 254.9975, 
    254.9969, 254.9973, 254.9972, 254.9975, 254.9996, 254.9991, 254.9996, 
    254.9996, 254.9996, 254.9999, 255.0001, 255.0005, 255.0004, 255.0001, 
    254.9995, 254.9997, 254.9992, 254.9993, 254.9987, 254.999, 254.9981, 
    254.9984, 254.9977, 254.9978, 254.9977, 254.9977, 254.9977, 254.9979, 
    254.9978, 254.998, 254.9989, 254.9986, 254.9995, 254.9999, 255.0003, 
    255.0006, 255.0005, 255.0005, 255.0001, 254.9998, 254.9996, 254.9994, 
    254.9993, 254.9988, 254.9986, 254.998, 254.9982, 254.998, 254.9979, 
    254.9976, 254.9977, 254.9976, 254.998, 254.9977, 254.9982, 254.9981, 
    254.9992, 254.9997, 254.9999, 255.0001, 255.0005, 255.0002, 255.0003, 
    255, 254.9998, 254.9999, 254.9994, 254.9996, 254.9985, 254.999, 254.9979, 
    254.9981, 254.9978, 254.998, 254.9977, 254.998, 254.9975, 254.9974, 
    254.9975, 254.9973, 254.998, 254.9977, 254.9999, 254.9999, 254.9999, 
    255.0002, 255.0002, 255.0005, 255.0002, 255.0001, 254.9998, 254.9997, 
    254.9995, 254.9992, 254.9989, 254.9984, 254.9981, 254.9979, 254.998, 
    254.9979, 254.998, 254.9981, 254.9975, 254.9978, 254.9973, 254.9973, 
    254.9976, 254.9973, 254.9999, 255, 255.0003, 255.0001, 255.0005, 
    255.0002, 255.0001, 254.9996, 254.9995, 254.9994, 254.9992, 254.9989, 
    254.9985, 254.9982, 254.9978, 254.9979, 254.9979, 254.9978, 254.998, 
    254.9978, 254.9977, 254.9978, 254.9973, 254.9975, 254.9973, 254.9974, 
    255, 254.9998, 254.9999, 254.9998, 254.9999, 254.9994, 254.9993, 
    254.9987, 254.9989, 254.9986, 254.9989, 254.9989, 254.9985, 254.9989, 
    254.9982, 254.9986, 254.9978, 254.9982, 254.9978, 254.9978, 254.9977, 
    254.9976, 254.9974, 254.9971, 254.9972, 254.997, 254.9996, 254.9994, 
    254.9995, 254.9993, 254.9991, 254.9989, 254.9984, 254.9986, 254.9983, 
    254.9982, 254.9987, 254.9984, 254.9993, 254.9992, 254.9993, 254.9996, 
    254.9985, 254.9991, 254.9981, 254.9984, 254.9976, 254.998, 254.9972, 
    254.9969, 254.9966, 254.9963, 254.9993, 254.9995, 254.9993, 254.999, 
    254.9987, 254.9984, 254.9984, 254.9983, 254.9981, 254.998, 254.9982, 
    254.998, 254.9991, 254.9985, 254.9995, 254.9992, 254.999, 254.9991, 
    254.9986, 254.9985, 254.998, 254.9983, 254.997, 254.9975, 254.9961, 
    254.9965, 254.9995, 254.9994, 254.9988, 254.9991, 254.9984, 254.9982, 
    254.998, 254.9979, 254.9978, 254.9978, 254.9979, 254.9978, 254.9984, 
    254.9981, 254.9989, 254.9987, 254.9988, 254.9989, 254.9986, 254.9982, 
    254.9983, 254.9981, 254.9978, 254.9984, 254.9969, 254.9977, 254.9992, 
    254.9989, 254.9988, 254.999, 254.9982, 254.9985, 254.9978, 254.9979, 
    254.9976, 254.9978, 254.9978, 254.998, 254.9981, 254.9985, 254.9987, 
    254.9989, 254.9989, 254.9986, 254.9982, 254.9978, 254.9979, 254.9977, 
    254.9984, 254.9981, 254.9982, 254.9979, 254.9986, 254.9979, 254.9987, 
    254.9987, 254.9985, 254.998, 254.998, 254.9979, 254.9979, 254.9982, 
    254.9983, 254.9985, 254.9985, 254.9987, 254.9988, 254.9987, 254.9986, 
    254.9982, 254.9979, 254.9976, 254.9975, 254.9971, 254.9974, 254.9969, 
    254.9973, 254.9966, 254.9979, 254.9973, 254.9985, 254.9984, 254.9981, 
    254.9976, 254.9979, 254.9976, 254.9983, 254.9986, 254.9987, 254.9989, 
    254.9987, 254.9988, 254.9986, 254.9986, 254.9982, 254.9984, 254.9978, 
    254.9976, 254.997, 254.9966, 254.9963, 254.9961, 254.9961, 254.9961 ;

 THBOT =
  256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044 ;

 TKE1 =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TLAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 TLAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TOTCOLC =
  18.24, 18.23998, 18.23999, 18.23998, 18.23998, 18.23997, 18.24, 18.23998, 
    18.23999, 18.24, 18.23996, 18.23998, 18.23993, 18.23995, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23988, 18.2399, 
    18.23987, 18.23989, 18.23988, 18.2399, 18.23997, 18.23996, 18.23997, 
    18.23997, 18.23997, 18.23998, 18.23999, 18.24, 18.24, 18.23999, 18.23997, 
    18.23998, 18.23996, 18.23996, 18.23994, 18.23995, 18.23992, 18.23993, 
    18.2399, 18.23991, 18.2399, 18.2399, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23995, 18.23994, 18.23997, 18.23998, 18.24, 18.24, 18.24, 
    18.24, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 18.23994, 
    18.23994, 18.23992, 18.23992, 18.23992, 18.23991, 18.2399, 18.2399, 
    18.2399, 18.23992, 18.2399, 18.23992, 18.23992, 18.23996, 18.23997, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23998, 18.23998, 
    18.23997, 18.23997, 18.23993, 18.23995, 18.23991, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.2399, 18.23989, 18.23989, 18.23989, 
    18.23991, 18.2399, 18.23998, 18.23998, 18.23998, 18.23999, 18.23999, 
    18.24, 18.23999, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 
    18.23995, 18.23993, 18.23992, 18.23991, 18.23992, 18.23991, 18.23992, 
    18.23992, 18.23989, 18.23991, 18.23989, 18.23989, 18.2399, 18.23989, 
    18.23998, 18.23998, 18.23999, 18.23999, 18.24, 18.23999, 18.23999, 
    18.23997, 18.23997, 18.23997, 18.23996, 18.23995, 18.23993, 18.23992, 
    18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.2399, 
    18.23991, 18.23989, 18.23989, 18.23989, 18.23989, 18.23998, 18.23998, 
    18.23998, 18.23998, 18.23998, 18.23997, 18.23996, 18.23994, 18.23995, 
    18.23994, 18.23995, 18.23995, 18.23994, 18.23995, 18.23992, 18.23994, 
    18.23991, 18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23989, 
    18.23988, 18.23988, 18.23987, 18.23997, 18.23997, 18.23997, 18.23996, 
    18.23996, 18.23995, 18.23993, 18.23994, 18.23993, 18.23992, 18.23994, 
    18.23993, 18.23996, 18.23996, 18.23996, 18.23997, 18.23993, 18.23995, 
    18.23992, 18.23993, 18.2399, 18.23991, 18.23989, 18.23987, 18.23986, 
    18.23985, 18.23996, 18.23997, 18.23996, 18.23995, 18.23994, 18.23993, 
    18.23993, 18.23993, 18.23992, 18.23991, 18.23993, 18.23991, 18.23996, 
    18.23993, 18.23997, 18.23996, 18.23995, 18.23995, 18.23994, 18.23993, 
    18.23992, 18.23993, 18.23988, 18.2399, 18.23984, 18.23985, 18.23997, 
    18.23996, 18.23994, 18.23995, 18.23993, 18.23992, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.23991, 18.23993, 18.23992, 18.23995, 
    18.23994, 18.23994, 18.23995, 18.23994, 18.23992, 18.23992, 18.23992, 
    18.23991, 18.23993, 18.23987, 18.23991, 18.23996, 18.23995, 18.23995, 
    18.23995, 18.23992, 18.23993, 18.23991, 18.23991, 18.2399, 18.23991, 
    18.23991, 18.23992, 18.23992, 18.23993, 18.23994, 18.23995, 18.23995, 
    18.23994, 18.23992, 18.23991, 18.23991, 18.2399, 18.23993, 18.23992, 
    18.23992, 18.23991, 18.23994, 18.23991, 18.23994, 18.23994, 18.23993, 
    18.23992, 18.23991, 18.23991, 18.23991, 18.23992, 18.23993, 18.23993, 
    18.23993, 18.23994, 18.23995, 18.23994, 18.23994, 18.23992, 18.23991, 
    18.2399, 18.23989, 18.23988, 18.23989, 18.23987, 18.23989, 18.23986, 
    18.23991, 18.23989, 18.23993, 18.23993, 18.23992, 18.2399, 18.23991, 
    18.2399, 18.23993, 18.23994, 18.23994, 18.23995, 18.23994, 18.23994, 
    18.23994, 18.23994, 18.23992, 18.23993, 18.23991, 18.2399, 18.23987, 
    18.23986, 18.23985, 18.23984, 18.23984, 18.23984 ;

 TOTCOLCH4 =
  1.38377e-05, 1.362747e-05, 1.366827e-05, 1.349928e-05, 1.359294e-05, 
    1.34824e-05, 1.379501e-05, 1.361914e-05, 1.373134e-05, 1.381875e-05, 
    1.317342e-05, 1.349176e-05, 1.284615e-05, 1.304669e-05, 1.263438e-05, 
    1.287725e-05, 1.256382e-05, 1.264453e-05, 1.240294e-05, 1.247176e-05, 
    1.216705e-05, 1.237129e-05, 1.201184e-05, 1.221556e-05, 1.218347e-05, 
    1.237808e-05, 1.342749e-05, 1.321289e-05, 1.344024e-05, 1.340955e-05, 
    1.342332e-05, 1.3591e-05, 1.367575e-05, 1.385382e-05, 1.382144e-05, 
    1.369069e-05, 1.339576e-05, 1.349564e-05, 1.324446e-05, 1.325012e-05, 
    1.297262e-05, 1.309743e-05, 1.272956e-05, 1.286921e-05, 1.246888e-05, 
    1.256862e-05, 1.247355e-05, 1.250231e-05, 1.247317e-05, 1.261971e-05, 
    1.255675e-05, 1.268633e-05, 1.307401e-05, 1.29322e-05, 1.335705e-05, 
    1.361501e-05, 1.378728e-05, 1.39099e-05, 1.389254e-05, 1.385948e-05, 
    1.368992e-05, 1.353111e-05, 1.34105e-05, 1.333003e-05, 1.325093e-05, 
    1.301259e-05, 1.288726e-05, 1.270145e-05, 1.275489e-05, 1.266447e-05, 
    1.257857e-05, 1.243541e-05, 1.245888e-05, 1.239614e-05, 1.266686e-05, 
    1.248639e-05, 1.278541e-05, 1.270307e-05, 1.322939e-05, 1.346867e-05, 
    1.357079e-05, 1.366042e-05, 1.38792e-05, 1.3728e-05, 1.378755e-05, 
    1.364603e-05, 1.355633e-05, 1.360067e-05, 1.332784e-05, 1.343368e-05, 
    1.287985e-05, 1.311721e-05, 1.258857e-05, 1.274391e-05, 1.255156e-05, 
    1.264943e-05, 1.248211e-05, 1.263261e-05, 1.237286e-05, 1.23169e-05, 
    1.235512e-05, 1.220891e-05, 1.2641e-05, 1.247354e-05, 1.360192e-05, 
    1.359468e-05, 1.3561e-05, 1.370926e-05, 1.371835e-05, 1.38547e-05, 
    1.373337e-05, 1.368179e-05, 1.355115e-05, 1.347406e-05, 1.340092e-05, 
    1.324063e-05, 1.306251e-05, 1.281524e-05, 1.273379e-05, 1.260858e-05, 
    1.268525e-05, 1.261754e-05, 1.269325e-05, 1.272885e-05, 1.233784e-05, 
    1.255616e-05, 1.222984e-05, 1.22477e-05, 1.239465e-05, 1.224569e-05, 
    1.35896e-05, 1.363125e-05, 1.377613e-05, 1.366271e-05, 1.386958e-05, 
    1.375366e-05, 1.368713e-05, 1.343145e-05, 1.337551e-05, 1.332369e-05, 
    1.32216e-05, 1.309103e-05, 1.286334e-05, 1.276346e-05, 1.257359e-05, 
    1.258743e-05, 1.258256e-05, 1.254042e-05, 1.2645e-05, 1.252332e-05, 
    1.250299e-05, 1.25562e-05, 1.22501e-05, 1.233688e-05, 1.224808e-05, 
    1.230452e-05, 1.361771e-05, 1.354768e-05, 1.35855e-05, 1.35144e-05, 
    1.356448e-05, 1.33423e-05, 1.327595e-05, 1.296726e-05, 1.309359e-05, 
    1.289281e-05, 1.307314e-05, 1.30411e-05, 1.288626e-05, 1.306337e-05, 
    1.277499e-05, 1.293851e-05, 1.253878e-05, 1.281418e-05, 1.252168e-05, 
    1.257441e-05, 1.248722e-05, 1.240955e-05, 1.231243e-05, 1.213502e-05, 
    1.217589e-05, 1.202891e-05, 1.344351e-05, 1.335311e-05, 1.336107e-05, 
    1.326669e-05, 1.319705e-05, 1.304664e-05, 1.280701e-05, 1.289688e-05, 
    1.283334e-05, 1.279809e-05, 1.294957e-05, 1.279554e-05, 1.329274e-05, 
    1.321185e-05, 1.325999e-05, 1.343637e-05, 1.287613e-05, 1.316241e-05, 
    1.273069e-05, 1.278946e-05, 1.242059e-05, 1.265462e-05, 1.219845e-05, 
    1.200795e-05, 1.183142e-05, 1.162854e-05, 1.330387e-05, 1.336519e-05, 
    1.325548e-05, 1.310426e-05, 1.296464e-05, 1.278007e-05, 1.286452e-05, 
    1.282768e-05, 1.273266e-05, 1.265317e-05, 1.281604e-05, 1.26333e-05, 
    1.319309e-05, 1.285142e-05, 1.33884e-05, 1.322573e-05, 1.311316e-05, 
    1.31625e-05, 1.290718e-05, 1.284733e-05, 1.269805e-05, 1.283131e-05, 
    1.205469e-05, 1.239318e-05, 1.147674e-05, 1.172545e-05, 1.338664e-05, 
    1.330409e-05, 1.301834e-05, 1.315398e-05, 1.287152e-05, 1.277072e-05, 
    1.268923e-05, 1.258563e-05, 1.257449e-05, 1.251348e-05, 1.261359e-05, 
    1.251743e-05, 1.277968e-05, 1.271931e-05, 1.305089e-05, 1.294671e-05, 
    1.299459e-05, 1.30472e-05, 1.288516e-05, 1.281346e-05, 1.280957e-05, 
    1.275103e-05, 1.258711e-05, 1.286985e-05, 1.201161e-05, 1.253571e-05, 
    1.321429e-05, 1.305625e-05, 1.303377e-05, 1.309485e-05, 1.27808e-05, 
    1.283151e-05, 1.251497e-05, 1.26287e-05, 1.244279e-05, 1.253489e-05, 
    1.254849e-05, 1.26677e-05, 1.274235e-05, 1.282468e-05, 1.297011e-05, 
    1.308598e-05, 1.3059e-05, 1.293186e-05, 1.280228e-05, 1.257348e-05, 
    1.262332e-05, 1.245684e-05, 1.279562e-05, 1.271346e-05, 1.278581e-05, 
    1.259781e-05, 1.289927e-05, 1.265867e-05, 1.298445e-05, 1.294774e-05, 
    1.283446e-05, 1.270078e-05, 1.264769e-05, 1.259117e-05, 1.262603e-05, 
    1.27961e-05, 1.282414e-05, 1.283722e-05, 1.286868e-05, 1.295573e-05, 
    1.302799e-05, 1.296196e-05, 1.289277e-05, 1.279604e-05, 1.260942e-05, 
    1.240844e-05, 1.235968e-05, 1.212914e-05, 1.231648e-05, 1.200874e-05, 
    1.226988e-05, 1.182132e-05, 1.263842e-05, 1.227768e-05, 1.282933e-05, 
    1.286508e-05, 1.273492e-05, 1.244031e-05, 1.259869e-05, 1.241364e-05, 
    1.282524e-05, 1.292748e-05, 1.298025e-05, 1.307892e-05, 1.297799e-05, 
    1.298619e-05, 1.288992e-05, 1.292082e-05, 1.278913e-05, 1.281411e-05, 
    1.254882e-05, 1.24151e-05, 1.204423e-05, 1.182217e-05, 1.160061e-05, 
    1.150429e-05, 1.147516e-05, 1.146301e-05 ;

 TOTCOLN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTECOSYSC =
  18.24, 18.23998, 18.23999, 18.23998, 18.23998, 18.23997, 18.24, 18.23998, 
    18.23999, 18.24, 18.23996, 18.23998, 18.23993, 18.23995, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23988, 18.2399, 
    18.23987, 18.23989, 18.23988, 18.2399, 18.23997, 18.23996, 18.23997, 
    18.23997, 18.23997, 18.23998, 18.23999, 18.24, 18.24, 18.23999, 18.23997, 
    18.23998, 18.23996, 18.23996, 18.23994, 18.23995, 18.23992, 18.23993, 
    18.2399, 18.23991, 18.2399, 18.2399, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23995, 18.23994, 18.23997, 18.23998, 18.24, 18.24, 18.24, 
    18.24, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 18.23994, 
    18.23994, 18.23992, 18.23992, 18.23992, 18.23991, 18.2399, 18.2399, 
    18.2399, 18.23992, 18.2399, 18.23992, 18.23992, 18.23996, 18.23997, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23998, 18.23998, 
    18.23997, 18.23997, 18.23993, 18.23995, 18.23991, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.2399, 18.23989, 18.23989, 18.23989, 
    18.23991, 18.2399, 18.23998, 18.23998, 18.23998, 18.23999, 18.23999, 
    18.24, 18.23999, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 
    18.23995, 18.23993, 18.23992, 18.23991, 18.23992, 18.23991, 18.23992, 
    18.23992, 18.23989, 18.23991, 18.23989, 18.23989, 18.2399, 18.23989, 
    18.23998, 18.23998, 18.23999, 18.23999, 18.24, 18.23999, 18.23999, 
    18.23997, 18.23997, 18.23997, 18.23996, 18.23995, 18.23993, 18.23992, 
    18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.2399, 
    18.23991, 18.23989, 18.23989, 18.23989, 18.23989, 18.23998, 18.23998, 
    18.23998, 18.23998, 18.23998, 18.23997, 18.23996, 18.23994, 18.23995, 
    18.23994, 18.23995, 18.23995, 18.23994, 18.23995, 18.23992, 18.23994, 
    18.23991, 18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23989, 
    18.23988, 18.23988, 18.23987, 18.23997, 18.23997, 18.23997, 18.23996, 
    18.23996, 18.23995, 18.23993, 18.23994, 18.23993, 18.23992, 18.23994, 
    18.23993, 18.23996, 18.23996, 18.23996, 18.23997, 18.23993, 18.23995, 
    18.23992, 18.23993, 18.2399, 18.23991, 18.23989, 18.23987, 18.23986, 
    18.23985, 18.23996, 18.23997, 18.23996, 18.23995, 18.23994, 18.23993, 
    18.23993, 18.23993, 18.23992, 18.23991, 18.23993, 18.23991, 18.23996, 
    18.23993, 18.23997, 18.23996, 18.23995, 18.23995, 18.23994, 18.23993, 
    18.23992, 18.23993, 18.23988, 18.2399, 18.23984, 18.23985, 18.23997, 
    18.23996, 18.23994, 18.23995, 18.23993, 18.23992, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.23991, 18.23993, 18.23992, 18.23995, 
    18.23994, 18.23994, 18.23995, 18.23994, 18.23992, 18.23992, 18.23992, 
    18.23991, 18.23993, 18.23987, 18.23991, 18.23996, 18.23995, 18.23995, 
    18.23995, 18.23992, 18.23993, 18.23991, 18.23991, 18.2399, 18.23991, 
    18.23991, 18.23992, 18.23992, 18.23993, 18.23994, 18.23995, 18.23995, 
    18.23994, 18.23992, 18.23991, 18.23991, 18.2399, 18.23993, 18.23992, 
    18.23992, 18.23991, 18.23994, 18.23991, 18.23994, 18.23994, 18.23993, 
    18.23992, 18.23991, 18.23991, 18.23991, 18.23992, 18.23993, 18.23993, 
    18.23993, 18.23994, 18.23995, 18.23994, 18.23994, 18.23992, 18.23991, 
    18.2399, 18.23989, 18.23988, 18.23989, 18.23987, 18.23989, 18.23986, 
    18.23991, 18.23989, 18.23993, 18.23993, 18.23992, 18.2399, 18.23991, 
    18.2399, 18.23993, 18.23994, 18.23994, 18.23995, 18.23994, 18.23994, 
    18.23994, 18.23994, 18.23992, 18.23993, 18.23991, 18.2399, 18.23987, 
    18.23986, 18.23985, 18.23984, 18.23984, 18.23984 ;

 TOTECOSYSN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTLITC =
  5.976202e-05, 5.976187e-05, 5.97619e-05, 5.976178e-05, 5.976185e-05, 
    5.976177e-05, 5.976199e-05, 5.976186e-05, 5.976194e-05, 5.9762e-05, 
    5.976155e-05, 5.976178e-05, 5.976132e-05, 5.976146e-05, 5.976111e-05, 
    5.976134e-05, 5.976106e-05, 5.976111e-05, 5.976095e-05, 5.9761e-05, 
    5.976079e-05, 5.976093e-05, 5.976068e-05, 5.976082e-05, 5.97608e-05, 
    5.976094e-05, 5.976173e-05, 5.976158e-05, 5.976174e-05, 5.976172e-05, 
    5.976173e-05, 5.976185e-05, 5.97619e-05, 5.976203e-05, 5.976201e-05, 
    5.976191e-05, 5.976171e-05, 5.976178e-05, 5.97616e-05, 5.976161e-05, 
    5.976141e-05, 5.97615e-05, 5.976117e-05, 5.976126e-05, 5.9761e-05, 
    5.976106e-05, 5.9761e-05, 5.976102e-05, 5.9761e-05, 5.97611e-05, 
    5.976106e-05, 5.976114e-05, 5.976148e-05, 5.976138e-05, 5.976168e-05, 
    5.976186e-05, 5.976198e-05, 5.976206e-05, 5.976205e-05, 5.976203e-05, 
    5.976191e-05, 5.97618e-05, 5.976172e-05, 5.976166e-05, 5.976161e-05, 
    5.976144e-05, 5.976135e-05, 5.976115e-05, 5.976119e-05, 5.976113e-05, 
    5.976107e-05, 5.976097e-05, 5.976099e-05, 5.976095e-05, 5.976113e-05, 
    5.976101e-05, 5.976121e-05, 5.976115e-05, 5.976159e-05, 5.976176e-05, 
    5.976183e-05, 5.976189e-05, 5.976205e-05, 5.976194e-05, 5.976198e-05, 
    5.976188e-05, 5.976182e-05, 5.976185e-05, 5.976166e-05, 5.976174e-05, 
    5.976135e-05, 5.976151e-05, 5.976108e-05, 5.976118e-05, 5.976105e-05, 
    5.976112e-05, 5.976101e-05, 5.976111e-05, 5.976093e-05, 5.976089e-05, 
    5.976092e-05, 5.976082e-05, 5.976111e-05, 5.9761e-05, 5.976185e-05, 
    5.976185e-05, 5.976182e-05, 5.976193e-05, 5.976193e-05, 5.976203e-05, 
    5.976194e-05, 5.976191e-05, 5.976182e-05, 5.976176e-05, 5.976171e-05, 
    5.97616e-05, 5.976147e-05, 5.97613e-05, 5.976118e-05, 5.976109e-05, 
    5.976114e-05, 5.97611e-05, 5.976115e-05, 5.976117e-05, 5.976091e-05, 
    5.976106e-05, 5.976083e-05, 5.976085e-05, 5.976095e-05, 5.976085e-05, 
    5.976184e-05, 5.976187e-05, 5.976197e-05, 5.976189e-05, 5.976204e-05, 
    5.976196e-05, 5.976191e-05, 5.976173e-05, 5.976169e-05, 5.976166e-05, 
    5.976159e-05, 5.97615e-05, 5.976133e-05, 5.976119e-05, 5.976107e-05, 
    5.976108e-05, 5.976107e-05, 5.976105e-05, 5.976111e-05, 5.976103e-05, 
    5.976102e-05, 5.976106e-05, 5.976085e-05, 5.976091e-05, 5.976085e-05, 
    5.976089e-05, 5.976186e-05, 5.976181e-05, 5.976184e-05, 5.976179e-05, 
    5.976183e-05, 5.976167e-05, 5.976162e-05, 5.976141e-05, 5.97615e-05, 
    5.976135e-05, 5.976148e-05, 5.976146e-05, 5.976135e-05, 5.976147e-05, 
    5.97612e-05, 5.976139e-05, 5.976105e-05, 5.976123e-05, 5.976103e-05, 
    5.976107e-05, 5.976101e-05, 5.976096e-05, 5.976089e-05, 5.976077e-05, 
    5.97608e-05, 5.976069e-05, 5.976174e-05, 5.976168e-05, 5.976169e-05, 
    5.976162e-05, 5.976157e-05, 5.976146e-05, 5.976129e-05, 5.976136e-05, 
    5.976124e-05, 5.976122e-05, 5.976139e-05, 5.976129e-05, 5.976163e-05, 
    5.976158e-05, 5.976161e-05, 5.976174e-05, 5.976134e-05, 5.976154e-05, 
    5.976117e-05, 5.976128e-05, 5.976097e-05, 5.976112e-05, 5.976081e-05, 
    5.976068e-05, 5.976055e-05, 5.976041e-05, 5.976165e-05, 5.976169e-05, 
    5.976161e-05, 5.97615e-05, 5.976141e-05, 5.976127e-05, 5.976126e-05, 
    5.976124e-05, 5.976117e-05, 5.976112e-05, 5.976123e-05, 5.976111e-05, 
    5.976157e-05, 5.976133e-05, 5.97617e-05, 5.976159e-05, 5.976151e-05, 
    5.976154e-05, 5.976137e-05, 5.976132e-05, 5.976115e-05, 5.976124e-05, 
    5.976071e-05, 5.976095e-05, 5.97603e-05, 5.976048e-05, 5.97617e-05, 
    5.976165e-05, 5.976145e-05, 5.976154e-05, 5.976127e-05, 5.97612e-05, 
    5.976114e-05, 5.976107e-05, 5.976107e-05, 5.976103e-05, 5.97611e-05, 
    5.976103e-05, 5.976127e-05, 5.976117e-05, 5.976147e-05, 5.976139e-05, 
    5.976143e-05, 5.976146e-05, 5.976135e-05, 5.976123e-05, 5.976123e-05, 
    5.976119e-05, 5.976108e-05, 5.976127e-05, 5.976068e-05, 5.976104e-05, 
    5.976158e-05, 5.976147e-05, 5.976146e-05, 5.97615e-05, 5.976121e-05, 
    5.976131e-05, 5.976103e-05, 5.97611e-05, 5.976098e-05, 5.976104e-05, 
    5.976105e-05, 5.976113e-05, 5.976118e-05, 5.976131e-05, 5.976141e-05, 
    5.976149e-05, 5.976147e-05, 5.976138e-05, 5.976122e-05, 5.976107e-05, 
    5.97611e-05, 5.976099e-05, 5.976129e-05, 5.976116e-05, 5.976121e-05, 
    5.976109e-05, 5.976136e-05, 5.976113e-05, 5.976142e-05, 5.976139e-05, 
    5.976131e-05, 5.976115e-05, 5.976112e-05, 5.976108e-05, 5.97611e-05, 
    5.976122e-05, 5.976123e-05, 5.976131e-05, 5.976134e-05, 5.97614e-05, 
    5.976145e-05, 5.976141e-05, 5.976135e-05, 5.976122e-05, 5.976109e-05, 
    5.976095e-05, 5.976092e-05, 5.976076e-05, 5.976089e-05, 5.976068e-05, 
    5.976086e-05, 5.976055e-05, 5.976111e-05, 5.976087e-05, 5.976131e-05, 
    5.976126e-05, 5.976118e-05, 5.976098e-05, 5.976109e-05, 5.976096e-05, 
    5.976123e-05, 5.976138e-05, 5.976142e-05, 5.976149e-05, 5.976142e-05, 
    5.976142e-05, 5.976135e-05, 5.976138e-05, 5.976121e-05, 5.97613e-05, 
    5.976105e-05, 5.976096e-05, 5.97607e-05, 5.976055e-05, 5.976039e-05, 
    5.976032e-05, 5.97603e-05, 5.976029e-05 ;

 TOTLITC_1m =
  5.976202e-05, 5.976187e-05, 5.97619e-05, 5.976178e-05, 5.976185e-05, 
    5.976177e-05, 5.976199e-05, 5.976186e-05, 5.976194e-05, 5.9762e-05, 
    5.976155e-05, 5.976178e-05, 5.976132e-05, 5.976146e-05, 5.976111e-05, 
    5.976134e-05, 5.976106e-05, 5.976111e-05, 5.976095e-05, 5.9761e-05, 
    5.976079e-05, 5.976093e-05, 5.976068e-05, 5.976082e-05, 5.97608e-05, 
    5.976094e-05, 5.976173e-05, 5.976158e-05, 5.976174e-05, 5.976172e-05, 
    5.976173e-05, 5.976185e-05, 5.97619e-05, 5.976203e-05, 5.976201e-05, 
    5.976191e-05, 5.976171e-05, 5.976178e-05, 5.97616e-05, 5.976161e-05, 
    5.976141e-05, 5.97615e-05, 5.976117e-05, 5.976126e-05, 5.9761e-05, 
    5.976106e-05, 5.9761e-05, 5.976102e-05, 5.9761e-05, 5.97611e-05, 
    5.976106e-05, 5.976114e-05, 5.976148e-05, 5.976138e-05, 5.976168e-05, 
    5.976186e-05, 5.976198e-05, 5.976206e-05, 5.976205e-05, 5.976203e-05, 
    5.976191e-05, 5.97618e-05, 5.976172e-05, 5.976166e-05, 5.976161e-05, 
    5.976144e-05, 5.976135e-05, 5.976115e-05, 5.976119e-05, 5.976113e-05, 
    5.976107e-05, 5.976097e-05, 5.976099e-05, 5.976095e-05, 5.976113e-05, 
    5.976101e-05, 5.976121e-05, 5.976115e-05, 5.976159e-05, 5.976176e-05, 
    5.976183e-05, 5.976189e-05, 5.976205e-05, 5.976194e-05, 5.976198e-05, 
    5.976188e-05, 5.976182e-05, 5.976185e-05, 5.976166e-05, 5.976174e-05, 
    5.976135e-05, 5.976151e-05, 5.976108e-05, 5.976118e-05, 5.976105e-05, 
    5.976112e-05, 5.976101e-05, 5.976111e-05, 5.976093e-05, 5.976089e-05, 
    5.976092e-05, 5.976082e-05, 5.976111e-05, 5.9761e-05, 5.976185e-05, 
    5.976185e-05, 5.976182e-05, 5.976193e-05, 5.976193e-05, 5.976203e-05, 
    5.976194e-05, 5.976191e-05, 5.976182e-05, 5.976176e-05, 5.976171e-05, 
    5.97616e-05, 5.976147e-05, 5.97613e-05, 5.976118e-05, 5.976109e-05, 
    5.976114e-05, 5.97611e-05, 5.976115e-05, 5.976117e-05, 5.976091e-05, 
    5.976106e-05, 5.976083e-05, 5.976085e-05, 5.976095e-05, 5.976085e-05, 
    5.976184e-05, 5.976187e-05, 5.976197e-05, 5.976189e-05, 5.976204e-05, 
    5.976196e-05, 5.976191e-05, 5.976173e-05, 5.976169e-05, 5.976166e-05, 
    5.976159e-05, 5.97615e-05, 5.976133e-05, 5.976119e-05, 5.976107e-05, 
    5.976108e-05, 5.976107e-05, 5.976105e-05, 5.976111e-05, 5.976103e-05, 
    5.976102e-05, 5.976106e-05, 5.976085e-05, 5.976091e-05, 5.976085e-05, 
    5.976089e-05, 5.976186e-05, 5.976181e-05, 5.976184e-05, 5.976179e-05, 
    5.976183e-05, 5.976167e-05, 5.976162e-05, 5.976141e-05, 5.97615e-05, 
    5.976135e-05, 5.976148e-05, 5.976146e-05, 5.976135e-05, 5.976147e-05, 
    5.97612e-05, 5.976139e-05, 5.976105e-05, 5.976123e-05, 5.976103e-05, 
    5.976107e-05, 5.976101e-05, 5.976096e-05, 5.976089e-05, 5.976077e-05, 
    5.97608e-05, 5.976069e-05, 5.976174e-05, 5.976168e-05, 5.976169e-05, 
    5.976162e-05, 5.976157e-05, 5.976146e-05, 5.976129e-05, 5.976136e-05, 
    5.976124e-05, 5.976122e-05, 5.976139e-05, 5.976129e-05, 5.976163e-05, 
    5.976158e-05, 5.976161e-05, 5.976174e-05, 5.976134e-05, 5.976154e-05, 
    5.976117e-05, 5.976128e-05, 5.976097e-05, 5.976112e-05, 5.976081e-05, 
    5.976068e-05, 5.976055e-05, 5.976041e-05, 5.976165e-05, 5.976169e-05, 
    5.976161e-05, 5.97615e-05, 5.976141e-05, 5.976127e-05, 5.976126e-05, 
    5.976124e-05, 5.976117e-05, 5.976112e-05, 5.976123e-05, 5.976111e-05, 
    5.976157e-05, 5.976133e-05, 5.97617e-05, 5.976159e-05, 5.976151e-05, 
    5.976154e-05, 5.976137e-05, 5.976132e-05, 5.976115e-05, 5.976124e-05, 
    5.976071e-05, 5.976095e-05, 5.97603e-05, 5.976048e-05, 5.97617e-05, 
    5.976165e-05, 5.976145e-05, 5.976154e-05, 5.976127e-05, 5.97612e-05, 
    5.976114e-05, 5.976107e-05, 5.976107e-05, 5.976103e-05, 5.97611e-05, 
    5.976103e-05, 5.976127e-05, 5.976117e-05, 5.976147e-05, 5.976139e-05, 
    5.976143e-05, 5.976146e-05, 5.976135e-05, 5.976123e-05, 5.976123e-05, 
    5.976119e-05, 5.976108e-05, 5.976127e-05, 5.976068e-05, 5.976104e-05, 
    5.976158e-05, 5.976147e-05, 5.976146e-05, 5.97615e-05, 5.976121e-05, 
    5.976131e-05, 5.976103e-05, 5.97611e-05, 5.976098e-05, 5.976104e-05, 
    5.976105e-05, 5.976113e-05, 5.976118e-05, 5.976131e-05, 5.976141e-05, 
    5.976149e-05, 5.976147e-05, 5.976138e-05, 5.976122e-05, 5.976107e-05, 
    5.97611e-05, 5.976099e-05, 5.976129e-05, 5.976116e-05, 5.976121e-05, 
    5.976109e-05, 5.976136e-05, 5.976113e-05, 5.976142e-05, 5.976139e-05, 
    5.976131e-05, 5.976115e-05, 5.976112e-05, 5.976108e-05, 5.97611e-05, 
    5.976122e-05, 5.976123e-05, 5.976131e-05, 5.976134e-05, 5.97614e-05, 
    5.976145e-05, 5.976141e-05, 5.976135e-05, 5.976122e-05, 5.976109e-05, 
    5.976095e-05, 5.976092e-05, 5.976076e-05, 5.976089e-05, 5.976068e-05, 
    5.976086e-05, 5.976055e-05, 5.976111e-05, 5.976087e-05, 5.976131e-05, 
    5.976126e-05, 5.976118e-05, 5.976098e-05, 5.976109e-05, 5.976096e-05, 
    5.976123e-05, 5.976138e-05, 5.976142e-05, 5.976149e-05, 5.976142e-05, 
    5.976142e-05, 5.976135e-05, 5.976138e-05, 5.976121e-05, 5.97613e-05, 
    5.976105e-05, 5.976096e-05, 5.97607e-05, 5.976055e-05, 5.976039e-05, 
    5.976032e-05, 5.97603e-05, 5.976029e-05 ;

 TOTLITN =
  1.375929e-06, 1.375925e-06, 1.375925e-06, 1.375922e-06, 1.375924e-06, 
    1.375922e-06, 1.375928e-06, 1.375924e-06, 1.375927e-06, 1.375928e-06, 
    1.375916e-06, 1.375922e-06, 1.375909e-06, 1.375913e-06, 1.375903e-06, 
    1.37591e-06, 1.375902e-06, 1.375903e-06, 1.375899e-06, 1.3759e-06, 
    1.375894e-06, 1.375898e-06, 1.375891e-06, 1.375895e-06, 1.375894e-06, 
    1.375898e-06, 1.375921e-06, 1.375916e-06, 1.375921e-06, 1.37592e-06, 
    1.375921e-06, 1.375924e-06, 1.375925e-06, 1.375929e-06, 1.375928e-06, 
    1.375926e-06, 1.37592e-06, 1.375922e-06, 1.375917e-06, 1.375917e-06, 
    1.375912e-06, 1.375914e-06, 1.375905e-06, 1.375907e-06, 1.3759e-06, 
    1.375902e-06, 1.3759e-06, 1.375901e-06, 1.3759e-06, 1.375903e-06, 
    1.375902e-06, 1.375904e-06, 1.375914e-06, 1.375911e-06, 1.375919e-06, 
    1.375924e-06, 1.375928e-06, 1.37593e-06, 1.37593e-06, 1.375929e-06, 
    1.375926e-06, 1.375923e-06, 1.37592e-06, 1.375919e-06, 1.375917e-06, 
    1.375912e-06, 1.37591e-06, 1.375904e-06, 1.375905e-06, 1.375904e-06, 
    1.375902e-06, 1.375899e-06, 1.3759e-06, 1.375899e-06, 1.375904e-06, 
    1.3759e-06, 1.375906e-06, 1.375904e-06, 1.375917e-06, 1.375921e-06, 
    1.375923e-06, 1.375925e-06, 1.375929e-06, 1.375926e-06, 1.375928e-06, 
    1.375925e-06, 1.375923e-06, 1.375924e-06, 1.375919e-06, 1.375921e-06, 
    1.37591e-06, 1.375915e-06, 1.375902e-06, 1.375905e-06, 1.375902e-06, 
    1.375903e-06, 1.3759e-06, 1.375903e-06, 1.375898e-06, 1.375897e-06, 
    1.375898e-06, 1.375895e-06, 1.375903e-06, 1.3759e-06, 1.375924e-06, 
    1.375924e-06, 1.375923e-06, 1.375926e-06, 1.375926e-06, 1.375929e-06, 
    1.375927e-06, 1.375926e-06, 1.375923e-06, 1.375921e-06, 1.37592e-06, 
    1.375917e-06, 1.375913e-06, 1.375908e-06, 1.375905e-06, 1.375903e-06, 
    1.375904e-06, 1.375903e-06, 1.375904e-06, 1.375905e-06, 1.375897e-06, 
    1.375902e-06, 1.375895e-06, 1.375896e-06, 1.375898e-06, 1.375896e-06, 
    1.375924e-06, 1.375925e-06, 1.375927e-06, 1.375925e-06, 1.375929e-06, 
    1.375927e-06, 1.375926e-06, 1.375921e-06, 1.37592e-06, 1.375918e-06, 
    1.375917e-06, 1.375914e-06, 1.375909e-06, 1.375906e-06, 1.375902e-06, 
    1.375902e-06, 1.375902e-06, 1.375901e-06, 1.375903e-06, 1.375901e-06, 
    1.375901e-06, 1.375902e-06, 1.375896e-06, 1.375897e-06, 1.375896e-06, 
    1.375897e-06, 1.375924e-06, 1.375923e-06, 1.375924e-06, 1.375922e-06, 
    1.375923e-06, 1.375919e-06, 1.375918e-06, 1.375912e-06, 1.375914e-06, 
    1.37591e-06, 1.375914e-06, 1.375913e-06, 1.37591e-06, 1.375913e-06, 
    1.375906e-06, 1.375911e-06, 1.375901e-06, 1.375906e-06, 1.375901e-06, 
    1.375902e-06, 1.3759e-06, 1.375899e-06, 1.375897e-06, 1.375893e-06, 
    1.375894e-06, 1.375891e-06, 1.375921e-06, 1.375919e-06, 1.375919e-06, 
    1.375917e-06, 1.375916e-06, 1.375913e-06, 1.375908e-06, 1.37591e-06, 
    1.375907e-06, 1.375906e-06, 1.375911e-06, 1.375908e-06, 1.375918e-06, 
    1.375916e-06, 1.375917e-06, 1.375921e-06, 1.37591e-06, 1.375915e-06, 
    1.375905e-06, 1.375908e-06, 1.375899e-06, 1.375903e-06, 1.375895e-06, 
    1.375891e-06, 1.375887e-06, 1.375883e-06, 1.375918e-06, 1.375919e-06, 
    1.375917e-06, 1.375914e-06, 1.375911e-06, 1.375908e-06, 1.375907e-06, 
    1.375907e-06, 1.375905e-06, 1.375903e-06, 1.375906e-06, 1.375903e-06, 
    1.375916e-06, 1.375909e-06, 1.37592e-06, 1.375917e-06, 1.375914e-06, 
    1.375915e-06, 1.37591e-06, 1.375909e-06, 1.375904e-06, 1.375907e-06, 
    1.375892e-06, 1.375898e-06, 1.37588e-06, 1.375885e-06, 1.37592e-06, 
    1.375918e-06, 1.375912e-06, 1.375915e-06, 1.375908e-06, 1.375906e-06, 
    1.375904e-06, 1.375902e-06, 1.375902e-06, 1.375901e-06, 1.375903e-06, 
    1.375901e-06, 1.375908e-06, 1.375905e-06, 1.375913e-06, 1.375911e-06, 
    1.375912e-06, 1.375913e-06, 1.37591e-06, 1.375906e-06, 1.375906e-06, 
    1.375905e-06, 1.375902e-06, 1.375907e-06, 1.375891e-06, 1.375901e-06, 
    1.375916e-06, 1.375913e-06, 1.375913e-06, 1.375914e-06, 1.375906e-06, 
    1.375909e-06, 1.375901e-06, 1.375903e-06, 1.375899e-06, 1.375901e-06, 
    1.375901e-06, 1.375904e-06, 1.375905e-06, 1.375909e-06, 1.375912e-06, 
    1.375914e-06, 1.375913e-06, 1.375911e-06, 1.375906e-06, 1.375902e-06, 
    1.375903e-06, 1.3759e-06, 1.375908e-06, 1.375905e-06, 1.375906e-06, 
    1.375902e-06, 1.37591e-06, 1.375903e-06, 1.375912e-06, 1.375911e-06, 
    1.375909e-06, 1.375904e-06, 1.375903e-06, 1.375902e-06, 1.375903e-06, 
    1.375906e-06, 1.375907e-06, 1.375909e-06, 1.37591e-06, 1.375911e-06, 
    1.375913e-06, 1.375911e-06, 1.37591e-06, 1.375906e-06, 1.375903e-06, 
    1.375899e-06, 1.375898e-06, 1.375893e-06, 1.375897e-06, 1.375891e-06, 
    1.375896e-06, 1.375887e-06, 1.375903e-06, 1.375896e-06, 1.375909e-06, 
    1.375907e-06, 1.375905e-06, 1.375899e-06, 1.375902e-06, 1.375899e-06, 
    1.375907e-06, 1.375911e-06, 1.375912e-06, 1.375914e-06, 1.375912e-06, 
    1.375912e-06, 1.37591e-06, 1.375911e-06, 1.375906e-06, 1.375908e-06, 
    1.375901e-06, 1.375899e-06, 1.375892e-06, 1.375887e-06, 1.375883e-06, 
    1.375881e-06, 1.37588e-06, 1.37588e-06 ;

 TOTLITN_1m =
  1.375929e-06, 1.375925e-06, 1.375925e-06, 1.375922e-06, 1.375924e-06, 
    1.375922e-06, 1.375928e-06, 1.375924e-06, 1.375927e-06, 1.375928e-06, 
    1.375916e-06, 1.375922e-06, 1.375909e-06, 1.375913e-06, 1.375903e-06, 
    1.37591e-06, 1.375902e-06, 1.375903e-06, 1.375899e-06, 1.3759e-06, 
    1.375894e-06, 1.375898e-06, 1.375891e-06, 1.375895e-06, 1.375894e-06, 
    1.375898e-06, 1.375921e-06, 1.375916e-06, 1.375921e-06, 1.37592e-06, 
    1.375921e-06, 1.375924e-06, 1.375925e-06, 1.375929e-06, 1.375928e-06, 
    1.375926e-06, 1.37592e-06, 1.375922e-06, 1.375917e-06, 1.375917e-06, 
    1.375912e-06, 1.375914e-06, 1.375905e-06, 1.375907e-06, 1.3759e-06, 
    1.375902e-06, 1.3759e-06, 1.375901e-06, 1.3759e-06, 1.375903e-06, 
    1.375902e-06, 1.375904e-06, 1.375914e-06, 1.375911e-06, 1.375919e-06, 
    1.375924e-06, 1.375928e-06, 1.37593e-06, 1.37593e-06, 1.375929e-06, 
    1.375926e-06, 1.375923e-06, 1.37592e-06, 1.375919e-06, 1.375917e-06, 
    1.375912e-06, 1.37591e-06, 1.375904e-06, 1.375905e-06, 1.375904e-06, 
    1.375902e-06, 1.375899e-06, 1.3759e-06, 1.375899e-06, 1.375904e-06, 
    1.3759e-06, 1.375906e-06, 1.375904e-06, 1.375917e-06, 1.375921e-06, 
    1.375923e-06, 1.375925e-06, 1.375929e-06, 1.375926e-06, 1.375928e-06, 
    1.375925e-06, 1.375923e-06, 1.375924e-06, 1.375919e-06, 1.375921e-06, 
    1.37591e-06, 1.375915e-06, 1.375902e-06, 1.375905e-06, 1.375902e-06, 
    1.375903e-06, 1.3759e-06, 1.375903e-06, 1.375898e-06, 1.375897e-06, 
    1.375898e-06, 1.375895e-06, 1.375903e-06, 1.3759e-06, 1.375924e-06, 
    1.375924e-06, 1.375923e-06, 1.375926e-06, 1.375926e-06, 1.375929e-06, 
    1.375927e-06, 1.375926e-06, 1.375923e-06, 1.375921e-06, 1.37592e-06, 
    1.375917e-06, 1.375913e-06, 1.375908e-06, 1.375905e-06, 1.375903e-06, 
    1.375904e-06, 1.375903e-06, 1.375904e-06, 1.375905e-06, 1.375897e-06, 
    1.375902e-06, 1.375895e-06, 1.375896e-06, 1.375898e-06, 1.375896e-06, 
    1.375924e-06, 1.375925e-06, 1.375927e-06, 1.375925e-06, 1.375929e-06, 
    1.375927e-06, 1.375926e-06, 1.375921e-06, 1.37592e-06, 1.375918e-06, 
    1.375917e-06, 1.375914e-06, 1.375909e-06, 1.375906e-06, 1.375902e-06, 
    1.375902e-06, 1.375902e-06, 1.375901e-06, 1.375903e-06, 1.375901e-06, 
    1.375901e-06, 1.375902e-06, 1.375896e-06, 1.375897e-06, 1.375896e-06, 
    1.375897e-06, 1.375924e-06, 1.375923e-06, 1.375924e-06, 1.375922e-06, 
    1.375923e-06, 1.375919e-06, 1.375918e-06, 1.375912e-06, 1.375914e-06, 
    1.37591e-06, 1.375914e-06, 1.375913e-06, 1.37591e-06, 1.375913e-06, 
    1.375906e-06, 1.375911e-06, 1.375901e-06, 1.375906e-06, 1.375901e-06, 
    1.375902e-06, 1.3759e-06, 1.375899e-06, 1.375897e-06, 1.375893e-06, 
    1.375894e-06, 1.375891e-06, 1.375921e-06, 1.375919e-06, 1.375919e-06, 
    1.375917e-06, 1.375916e-06, 1.375913e-06, 1.375908e-06, 1.37591e-06, 
    1.375907e-06, 1.375906e-06, 1.375911e-06, 1.375908e-06, 1.375918e-06, 
    1.375916e-06, 1.375917e-06, 1.375921e-06, 1.37591e-06, 1.375915e-06, 
    1.375905e-06, 1.375908e-06, 1.375899e-06, 1.375903e-06, 1.375895e-06, 
    1.375891e-06, 1.375887e-06, 1.375883e-06, 1.375918e-06, 1.375919e-06, 
    1.375917e-06, 1.375914e-06, 1.375911e-06, 1.375908e-06, 1.375907e-06, 
    1.375907e-06, 1.375905e-06, 1.375903e-06, 1.375906e-06, 1.375903e-06, 
    1.375916e-06, 1.375909e-06, 1.37592e-06, 1.375917e-06, 1.375914e-06, 
    1.375915e-06, 1.37591e-06, 1.375909e-06, 1.375904e-06, 1.375907e-06, 
    1.375892e-06, 1.375898e-06, 1.37588e-06, 1.375885e-06, 1.37592e-06, 
    1.375918e-06, 1.375912e-06, 1.375915e-06, 1.375908e-06, 1.375906e-06, 
    1.375904e-06, 1.375902e-06, 1.375902e-06, 1.375901e-06, 1.375903e-06, 
    1.375901e-06, 1.375908e-06, 1.375905e-06, 1.375913e-06, 1.375911e-06, 
    1.375912e-06, 1.375913e-06, 1.37591e-06, 1.375906e-06, 1.375906e-06, 
    1.375905e-06, 1.375902e-06, 1.375907e-06, 1.375891e-06, 1.375901e-06, 
    1.375916e-06, 1.375913e-06, 1.375913e-06, 1.375914e-06, 1.375906e-06, 
    1.375909e-06, 1.375901e-06, 1.375903e-06, 1.375899e-06, 1.375901e-06, 
    1.375901e-06, 1.375904e-06, 1.375905e-06, 1.375909e-06, 1.375912e-06, 
    1.375914e-06, 1.375913e-06, 1.375911e-06, 1.375906e-06, 1.375902e-06, 
    1.375903e-06, 1.3759e-06, 1.375908e-06, 1.375905e-06, 1.375906e-06, 
    1.375902e-06, 1.37591e-06, 1.375903e-06, 1.375912e-06, 1.375911e-06, 
    1.375909e-06, 1.375904e-06, 1.375903e-06, 1.375902e-06, 1.375903e-06, 
    1.375906e-06, 1.375907e-06, 1.375909e-06, 1.37591e-06, 1.375911e-06, 
    1.375913e-06, 1.375911e-06, 1.37591e-06, 1.375906e-06, 1.375903e-06, 
    1.375899e-06, 1.375898e-06, 1.375893e-06, 1.375897e-06, 1.375891e-06, 
    1.375896e-06, 1.375887e-06, 1.375903e-06, 1.375896e-06, 1.375909e-06, 
    1.375907e-06, 1.375905e-06, 1.375899e-06, 1.375902e-06, 1.375899e-06, 
    1.375907e-06, 1.375911e-06, 1.375912e-06, 1.375914e-06, 1.375912e-06, 
    1.375912e-06, 1.37591e-06, 1.375911e-06, 1.375906e-06, 1.375908e-06, 
    1.375901e-06, 1.375899e-06, 1.375892e-06, 1.375887e-06, 1.375883e-06, 
    1.375881e-06, 1.37588e-06, 1.37588e-06 ;

 TOTPFTC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTPFTN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TOTPRODC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTPRODN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTSOMC =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34457, 17.34459, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.3446, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34456, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34452, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.3445, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.34449, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34457, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34453, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34456, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34455, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 TOTSOMC_1m =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34457, 17.34459, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.3446, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34456, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34452, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.3445, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.34449, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34457, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34453, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34456, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34455, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 TOTSOMN =
  1.773759, 1.773758, 1.773758, 1.773756, 1.773757, 1.773756, 1.773759, 
    1.773757, 1.773759, 1.773759, 1.773753, 1.773756, 1.77375, 1.773752, 
    1.773747, 1.773751, 1.773747, 1.773747, 1.773745, 1.773746, 1.773743, 
    1.773745, 1.773742, 1.773744, 1.773743, 1.773745, 1.773756, 1.773754, 
    1.773756, 1.773756, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773758, 1.773755, 1.773756, 1.773754, 1.773754, 1.773751, 1.773753, 
    1.773748, 1.773749, 1.773746, 1.773747, 1.773746, 1.773746, 1.773746, 
    1.773747, 1.773747, 1.773748, 1.773752, 1.773751, 1.773755, 1.773757, 
    1.773759, 1.77376, 1.77376, 1.77376, 1.773758, 1.773757, 1.773756, 
    1.773755, 1.773754, 1.773752, 1.773751, 1.773748, 1.773749, 1.773748, 
    1.773747, 1.773746, 1.773746, 1.773745, 1.773748, 1.773746, 1.773749, 
    1.773748, 1.773754, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773759, 1.773758, 1.773757, 1.773757, 1.773755, 1.773756, 1.773751, 
    1.773753, 1.773747, 1.773748, 1.773747, 1.773748, 1.773746, 1.773747, 
    1.773745, 1.773744, 1.773745, 1.773744, 1.773747, 1.773746, 1.773757, 
    1.773757, 1.773757, 1.773758, 1.773758, 1.77376, 1.773759, 1.773758, 
    1.773757, 1.773756, 1.773755, 1.773754, 1.773752, 1.77375, 1.773748, 
    1.773747, 1.773748, 1.773747, 1.773748, 1.773748, 1.773745, 1.773747, 
    1.773744, 1.773744, 1.773745, 1.773744, 1.773757, 1.773758, 1.773759, 
    1.773758, 1.77376, 1.773759, 1.773758, 1.773756, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.77375, 1.773749, 1.773747, 1.773747, 1.773747, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773744, 1.773745, 
    1.773744, 1.773744, 1.773757, 1.773757, 1.773757, 1.773757, 1.773757, 
    1.773755, 1.773754, 1.773751, 1.773753, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773752, 1.773749, 1.773751, 1.773746, 1.773749, 1.773746, 
    1.773747, 1.773746, 1.773745, 1.773744, 1.773743, 1.773743, 1.773742, 
    1.773756, 1.773755, 1.773755, 1.773754, 1.773754, 1.773752, 1.77375, 
    1.773751, 1.773749, 1.773749, 1.773751, 1.77375, 1.773754, 1.773754, 
    1.773754, 1.773756, 1.773751, 1.773753, 1.773748, 1.77375, 1.773745, 
    1.773748, 1.773743, 1.773742, 1.77374, 1.773738, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.773751, 1.77375, 1.773749, 1.773749, 1.773748, 
    1.773748, 1.773749, 1.773747, 1.773754, 1.77375, 1.773755, 1.773754, 
    1.773753, 1.773753, 1.773751, 1.77375, 1.773748, 1.773749, 1.773742, 
    1.773745, 1.773736, 1.773739, 1.773755, 1.773755, 1.773752, 1.773753, 
    1.773749, 1.773749, 1.773748, 1.773747, 1.773747, 1.773746, 1.773747, 
    1.773746, 1.77375, 1.773748, 1.773752, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773749, 1.773749, 1.773748, 1.773747, 1.773749, 1.773742, 
    1.773746, 1.773754, 1.773752, 1.773752, 1.773753, 1.773749, 1.77375, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773748, 1.773748, 
    1.77375, 1.773751, 1.773752, 1.773752, 1.773751, 1.773749, 1.773747, 
    1.773747, 1.773746, 1.77375, 1.773748, 1.773749, 1.773747, 1.773751, 
    1.773748, 1.773751, 1.773751, 1.77375, 1.773748, 1.773747, 1.773747, 
    1.773747, 1.773749, 1.773749, 1.77375, 1.77375, 1.773751, 1.773752, 
    1.773751, 1.773751, 1.773749, 1.773747, 1.773745, 1.773745, 1.773743, 
    1.773744, 1.773742, 1.773744, 1.77374, 1.773747, 1.773744, 1.77375, 
    1.773749, 1.773748, 1.773746, 1.773747, 1.773745, 1.773749, 1.773751, 
    1.773751, 1.773752, 1.773751, 1.773752, 1.773751, 1.773751, 1.773749, 
    1.77375, 1.773747, 1.773745, 1.773742, 1.77374, 1.773738, 1.773737, 
    1.773736, 1.773736 ;

 TOTSOMN_1m =
  1.773759, 1.773758, 1.773758, 1.773756, 1.773757, 1.773756, 1.773759, 
    1.773757, 1.773759, 1.773759, 1.773753, 1.773756, 1.77375, 1.773752, 
    1.773747, 1.773751, 1.773747, 1.773747, 1.773745, 1.773746, 1.773743, 
    1.773745, 1.773742, 1.773744, 1.773743, 1.773745, 1.773756, 1.773754, 
    1.773756, 1.773756, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773758, 1.773755, 1.773756, 1.773754, 1.773754, 1.773751, 1.773753, 
    1.773748, 1.773749, 1.773746, 1.773747, 1.773746, 1.773746, 1.773746, 
    1.773747, 1.773747, 1.773748, 1.773752, 1.773751, 1.773755, 1.773757, 
    1.773759, 1.77376, 1.77376, 1.77376, 1.773758, 1.773757, 1.773756, 
    1.773755, 1.773754, 1.773752, 1.773751, 1.773748, 1.773749, 1.773748, 
    1.773747, 1.773746, 1.773746, 1.773745, 1.773748, 1.773746, 1.773749, 
    1.773748, 1.773754, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773759, 1.773758, 1.773757, 1.773757, 1.773755, 1.773756, 1.773751, 
    1.773753, 1.773747, 1.773748, 1.773747, 1.773748, 1.773746, 1.773747, 
    1.773745, 1.773744, 1.773745, 1.773744, 1.773747, 1.773746, 1.773757, 
    1.773757, 1.773757, 1.773758, 1.773758, 1.77376, 1.773759, 1.773758, 
    1.773757, 1.773756, 1.773755, 1.773754, 1.773752, 1.77375, 1.773748, 
    1.773747, 1.773748, 1.773747, 1.773748, 1.773748, 1.773745, 1.773747, 
    1.773744, 1.773744, 1.773745, 1.773744, 1.773757, 1.773758, 1.773759, 
    1.773758, 1.77376, 1.773759, 1.773758, 1.773756, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.77375, 1.773749, 1.773747, 1.773747, 1.773747, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773744, 1.773745, 
    1.773744, 1.773744, 1.773757, 1.773757, 1.773757, 1.773757, 1.773757, 
    1.773755, 1.773754, 1.773751, 1.773753, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773752, 1.773749, 1.773751, 1.773746, 1.773749, 1.773746, 
    1.773747, 1.773746, 1.773745, 1.773744, 1.773743, 1.773743, 1.773742, 
    1.773756, 1.773755, 1.773755, 1.773754, 1.773754, 1.773752, 1.77375, 
    1.773751, 1.773749, 1.773749, 1.773751, 1.77375, 1.773754, 1.773754, 
    1.773754, 1.773756, 1.773751, 1.773753, 1.773748, 1.77375, 1.773745, 
    1.773748, 1.773743, 1.773742, 1.77374, 1.773738, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.773751, 1.77375, 1.773749, 1.773749, 1.773748, 
    1.773748, 1.773749, 1.773747, 1.773754, 1.77375, 1.773755, 1.773754, 
    1.773753, 1.773753, 1.773751, 1.77375, 1.773748, 1.773749, 1.773742, 
    1.773745, 1.773736, 1.773739, 1.773755, 1.773755, 1.773752, 1.773753, 
    1.773749, 1.773749, 1.773748, 1.773747, 1.773747, 1.773746, 1.773747, 
    1.773746, 1.77375, 1.773748, 1.773752, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773749, 1.773749, 1.773748, 1.773747, 1.773749, 1.773742, 
    1.773746, 1.773754, 1.773752, 1.773752, 1.773753, 1.773749, 1.77375, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773748, 1.773748, 
    1.77375, 1.773751, 1.773752, 1.773752, 1.773751, 1.773749, 1.773747, 
    1.773747, 1.773746, 1.77375, 1.773748, 1.773749, 1.773747, 1.773751, 
    1.773748, 1.773751, 1.773751, 1.77375, 1.773748, 1.773747, 1.773747, 
    1.773747, 1.773749, 1.773749, 1.77375, 1.77375, 1.773751, 1.773752, 
    1.773751, 1.773751, 1.773749, 1.773747, 1.773745, 1.773745, 1.773743, 
    1.773744, 1.773742, 1.773744, 1.77374, 1.773747, 1.773744, 1.77375, 
    1.773749, 1.773748, 1.773746, 1.773747, 1.773745, 1.773749, 1.773751, 
    1.773751, 1.773752, 1.773751, 1.773752, 1.773751, 1.773751, 1.773749, 
    1.77375, 1.773747, 1.773745, 1.773742, 1.77374, 1.773738, 1.773737, 
    1.773736, 1.773736 ;

 TOTVEGC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTVEGN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TREFMNAV =
  243.0876, 243.0908, 243.0902, 243.0928, 243.0914, 243.093, 243.0883, 
    243.0909, 243.0892, 243.0879, 243.0977, 243.0929, 243.1028, 243.0998, 
    243.1075, 243.1023, 243.1086, 243.1074, 243.111, 243.11, 243.1144, 
    243.1115, 243.1168, 243.1138, 243.1142, 243.1114, 243.0939, 243.0971, 
    243.0937, 243.0942, 243.094, 243.0914, 243.09, 243.0874, 243.0879, 
    243.0898, 243.0944, 243.0929, 243.0968, 243.0967, 243.1009, 243.099, 
    243.1062, 243.1042, 243.11, 243.1085, 243.1099, 243.1095, 243.11, 
    243.1078, 243.1087, 243.1068, 243.0994, 243.1015, 243.095, 243.0909, 
    243.0884, 243.0865, 243.0868, 243.0873, 243.0899, 243.0923, 243.0942, 
    243.0954, 243.0966, 243.1002, 243.1022, 243.1066, 243.1058, 243.1071, 
    243.1084, 243.1105, 243.1102, 243.1111, 243.1071, 243.1097, 243.1054, 
    243.1066, 243.0968, 243.0933, 243.0916, 243.0903, 243.087, 243.0893, 
    243.0884, 243.0906, 243.0919, 243.0913, 243.0955, 243.0938, 243.1023, 
    243.0987, 243.1082, 243.106, 243.1088, 243.1074, 243.1098, 243.1076, 
    243.1114, 243.1122, 243.1117, 243.1139, 243.1075, 243.1099, 243.0912, 
    243.0914, 243.0919, 243.0896, 243.0894, 243.0874, 243.0892, 243.09, 
    243.092, 243.0932, 243.0943, 243.0968, 243.0995, 243.1033, 243.1061, 
    243.108, 243.1068, 243.1078, 243.1067, 243.1062, 243.1119, 243.1087, 
    243.1136, 243.1133, 243.1111, 243.1133, 243.0914, 243.0908, 243.0885, 
    243.0903, 243.0871, 243.0889, 243.0899, 243.0938, 243.0947, 243.0955, 
    243.0971, 243.0991, 243.1026, 243.1057, 243.1085, 243.1083, 243.1084, 
    243.109, 243.1074, 243.1092, 243.1095, 243.1087, 243.1133, 243.112, 
    243.1133, 243.1125, 243.091, 243.0921, 243.0915, 243.0926, 243.0918, 
    243.0952, 243.0962, 243.101, 243.0991, 243.1021, 243.0994, 243.0999, 
    243.1022, 243.0995, 243.1055, 243.1014, 243.109, 243.1049, 243.1092, 
    243.1085, 243.1098, 243.1109, 243.1123, 243.115, 243.1144, 243.1166, 
    243.0937, 243.095, 243.095, 243.0964, 243.0975, 243.0998, 243.1035, 
    243.1021, 243.1047, 243.1052, 243.1013, 243.1037, 243.096, 243.0972, 
    243.0965, 243.0938, 243.1024, 243.098, 243.1062, 243.1038, 243.1107, 
    243.1072, 243.114, 243.1168, 243.1196, 243.1227, 243.0958, 243.0949, 
    243.0966, 243.0989, 243.1011, 243.1039, 243.1042, 243.1048, 243.1062, 
    243.1073, 243.1049, 243.1076, 243.0974, 243.1028, 243.0945, 243.097, 
    243.0987, 243.098, 243.102, 243.1029, 243.1066, 243.1047, 243.1161, 
    243.1111, 243.1251, 243.1212, 243.0946, 243.0958, 243.1002, 243.0981, 
    243.1041, 243.1056, 243.1068, 243.1083, 243.1085, 243.1093, 243.1079, 
    243.1093, 243.1039, 243.1063, 243.0997, 243.1013, 243.1006, 243.0998, 
    243.1023, 243.1049, 243.105, 243.1059, 243.1081, 243.1042, 243.1166, 
    243.1089, 243.0972, 243.0996, 243.1, 243.0991, 243.1054, 243.1031, 
    243.1093, 243.1077, 243.1104, 243.109, 243.1088, 243.1071, 243.106, 
    243.1032, 243.101, 243.0992, 243.0996, 243.1015, 243.1051, 243.1085, 
    243.1077, 243.1102, 243.1037, 243.1064, 243.1053, 243.1081, 243.1021, 
    243.1071, 243.1008, 243.1013, 243.1031, 243.1065, 243.1074, 243.1082, 
    243.1077, 243.1052, 243.1048, 243.103, 243.1025, 243.1012, 243.1001, 
    243.1011, 243.1022, 243.1052, 243.1079, 243.1109, 243.1116, 243.1149, 
    243.1122, 243.1167, 243.1127, 243.1196, 243.1074, 243.1127, 243.1032, 
    243.1042, 243.1061, 243.1104, 243.1081, 243.1108, 243.1048, 243.1016, 
    243.1008, 243.0993, 243.1009, 243.1007, 243.1022, 243.1018, 243.1053, 
    243.1034, 243.1088, 243.1108, 243.1163, 243.1197, 243.1232, 243.1247, 
    243.1251, 243.1253 ;

 TREFMNAV_R =
  243.0876, 243.0908, 243.0902, 243.0928, 243.0914, 243.093, 243.0883, 
    243.0909, 243.0892, 243.0879, 243.0977, 243.0929, 243.1028, 243.0998, 
    243.1075, 243.1023, 243.1086, 243.1074, 243.111, 243.11, 243.1144, 
    243.1115, 243.1168, 243.1138, 243.1142, 243.1114, 243.0939, 243.0971, 
    243.0937, 243.0942, 243.094, 243.0914, 243.09, 243.0874, 243.0879, 
    243.0898, 243.0944, 243.0929, 243.0968, 243.0967, 243.1009, 243.099, 
    243.1062, 243.1042, 243.11, 243.1085, 243.1099, 243.1095, 243.11, 
    243.1078, 243.1087, 243.1068, 243.0994, 243.1015, 243.095, 243.0909, 
    243.0884, 243.0865, 243.0868, 243.0873, 243.0899, 243.0923, 243.0942, 
    243.0954, 243.0966, 243.1002, 243.1022, 243.1066, 243.1058, 243.1071, 
    243.1084, 243.1105, 243.1102, 243.1111, 243.1071, 243.1097, 243.1054, 
    243.1066, 243.0968, 243.0933, 243.0916, 243.0903, 243.087, 243.0893, 
    243.0884, 243.0906, 243.0919, 243.0913, 243.0955, 243.0938, 243.1023, 
    243.0987, 243.1082, 243.106, 243.1088, 243.1074, 243.1098, 243.1076, 
    243.1114, 243.1122, 243.1117, 243.1139, 243.1075, 243.1099, 243.0912, 
    243.0914, 243.0919, 243.0896, 243.0894, 243.0874, 243.0892, 243.09, 
    243.092, 243.0932, 243.0943, 243.0968, 243.0995, 243.1033, 243.1061, 
    243.108, 243.1068, 243.1078, 243.1067, 243.1062, 243.1119, 243.1087, 
    243.1136, 243.1133, 243.1111, 243.1133, 243.0914, 243.0908, 243.0885, 
    243.0903, 243.0871, 243.0889, 243.0899, 243.0938, 243.0947, 243.0955, 
    243.0971, 243.0991, 243.1026, 243.1057, 243.1085, 243.1083, 243.1084, 
    243.109, 243.1074, 243.1092, 243.1095, 243.1087, 243.1133, 243.112, 
    243.1133, 243.1125, 243.091, 243.0921, 243.0915, 243.0926, 243.0918, 
    243.0952, 243.0962, 243.101, 243.0991, 243.1021, 243.0994, 243.0999, 
    243.1022, 243.0995, 243.1055, 243.1014, 243.109, 243.1049, 243.1092, 
    243.1085, 243.1098, 243.1109, 243.1123, 243.115, 243.1144, 243.1166, 
    243.0937, 243.095, 243.095, 243.0964, 243.0975, 243.0998, 243.1035, 
    243.1021, 243.1047, 243.1052, 243.1013, 243.1037, 243.096, 243.0972, 
    243.0965, 243.0938, 243.1024, 243.098, 243.1062, 243.1038, 243.1107, 
    243.1072, 243.114, 243.1168, 243.1196, 243.1227, 243.0958, 243.0949, 
    243.0966, 243.0989, 243.1011, 243.1039, 243.1042, 243.1048, 243.1062, 
    243.1073, 243.1049, 243.1076, 243.0974, 243.1028, 243.0945, 243.097, 
    243.0987, 243.098, 243.102, 243.1029, 243.1066, 243.1047, 243.1161, 
    243.1111, 243.1251, 243.1212, 243.0946, 243.0958, 243.1002, 243.0981, 
    243.1041, 243.1056, 243.1068, 243.1083, 243.1085, 243.1093, 243.1079, 
    243.1093, 243.1039, 243.1063, 243.0997, 243.1013, 243.1006, 243.0998, 
    243.1023, 243.1049, 243.105, 243.1059, 243.1081, 243.1042, 243.1166, 
    243.1089, 243.0972, 243.0996, 243.1, 243.0991, 243.1054, 243.1031, 
    243.1093, 243.1077, 243.1104, 243.109, 243.1088, 243.1071, 243.106, 
    243.1032, 243.101, 243.0992, 243.0996, 243.1015, 243.1051, 243.1085, 
    243.1077, 243.1102, 243.1037, 243.1064, 243.1053, 243.1081, 243.1021, 
    243.1071, 243.1008, 243.1013, 243.1031, 243.1065, 243.1074, 243.1082, 
    243.1077, 243.1052, 243.1048, 243.103, 243.1025, 243.1012, 243.1001, 
    243.1011, 243.1022, 243.1052, 243.1079, 243.1109, 243.1116, 243.1149, 
    243.1122, 243.1167, 243.1127, 243.1196, 243.1074, 243.1127, 243.1032, 
    243.1042, 243.1061, 243.1104, 243.1081, 243.1108, 243.1048, 243.1016, 
    243.1008, 243.0993, 243.1009, 243.1007, 243.1022, 243.1018, 243.1053, 
    243.1034, 243.1088, 243.1108, 243.1163, 243.1197, 243.1232, 243.1247, 
    243.1251, 243.1253 ;

 TREFMNAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TREFMXAV =
  270.7643, 270.7622, 270.7626, 270.7609, 270.7618, 270.7607, 270.7638, 
    270.7621, 270.7632, 270.7641, 270.7577, 270.7608, 270.7543, 270.7563, 
    270.7512, 270.7546, 270.7505, 270.7512, 270.7488, 270.7495, 270.7466, 
    270.7485, 270.745, 270.747, 270.7467, 270.7486, 270.7601, 270.7581, 
    270.7603, 270.76, 270.7601, 270.7618, 270.7627, 270.7644, 270.7641, 
    270.7628, 270.7598, 270.7608, 270.7583, 270.7583, 270.7555, 270.7568, 
    270.752, 270.7534, 270.7495, 270.7505, 270.7495, 270.7498, 270.7495, 
    270.751, 270.7504, 270.7516, 270.7566, 270.7551, 270.7594, 270.7621, 
    270.7638, 270.765, 270.7648, 270.7645, 270.7628, 270.7612, 270.7599, 
    270.7592, 270.7583, 270.756, 270.7547, 270.7518, 270.7523, 270.7514, 
    270.7506, 270.7492, 270.7494, 270.7488, 270.7514, 270.7497, 270.7526, 
    270.7518, 270.7583, 270.7606, 270.7617, 270.7625, 270.7647, 270.7632, 
    270.7638, 270.7623, 270.7614, 270.7619, 270.7591, 270.7602, 270.7546, 
    270.757, 270.7507, 270.7522, 270.7503, 270.7513, 270.7496, 270.7511, 
    270.7485, 270.748, 270.7484, 270.7469, 270.7512, 270.7495, 270.7619, 
    270.7618, 270.7615, 270.763, 270.7631, 270.7644, 270.7632, 270.7627, 
    270.7614, 270.7606, 270.7599, 270.7582, 270.7565, 270.7539, 270.7521, 
    270.7509, 270.7516, 270.7509, 270.7517, 270.752, 270.7482, 270.7504, 
    270.7471, 270.7473, 270.7488, 270.7473, 270.7618, 270.7622, 270.7636, 
    270.7625, 270.7646, 270.7634, 270.7628, 270.7602, 270.7596, 270.7591, 
    270.7581, 270.7567, 270.7544, 270.7524, 270.7505, 270.7506, 270.7506, 
    270.7502, 270.7512, 270.75, 270.7498, 270.7504, 270.7473, 270.7482, 
    270.7473, 270.7479, 270.7621, 270.7614, 270.7617, 270.761, 270.7615, 
    270.7593, 270.7586, 270.7555, 270.7568, 270.7547, 270.7565, 270.7562, 
    270.7547, 270.7564, 270.7525, 270.7552, 270.7502, 270.7529, 270.75, 
    270.7505, 270.7497, 270.7489, 270.748, 270.7462, 270.7466, 270.7451, 
    270.7603, 270.7594, 270.7595, 270.7585, 270.7578, 270.7563, 270.7538, 
    270.7547, 270.7531, 270.7527, 270.7553, 270.7537, 270.7588, 270.758, 
    270.7585, 270.7602, 270.7546, 270.7575, 270.7521, 270.7536, 270.749, 
    270.7513, 270.7468, 270.7449, 270.7431, 270.741, 270.7589, 270.7595, 
    270.7584, 270.7569, 270.7554, 270.7535, 270.7533, 270.753, 270.7521, 
    270.7513, 270.7529, 270.7511, 270.7579, 270.7543, 270.7597, 270.7581, 
    270.757, 270.7574, 270.7548, 270.7542, 270.7518, 270.753, 270.7454, 
    270.7488, 270.7394, 270.742, 270.7597, 270.7589, 270.756, 270.7574, 
    270.7534, 270.7524, 270.7516, 270.7506, 270.7505, 270.7499, 270.7509, 
    270.75, 270.7535, 270.752, 270.7563, 270.7552, 270.7557, 270.7563, 
    270.7546, 270.7529, 270.7528, 270.7523, 270.7508, 270.7534, 270.7451, 
    270.7503, 270.758, 270.7564, 270.7561, 270.7567, 270.7525, 270.7541, 
    270.7499, 270.7511, 270.7492, 270.7502, 270.7503, 270.7514, 270.7522, 
    270.754, 270.7555, 270.7567, 270.7564, 270.7551, 270.7528, 270.7505, 
    270.751, 270.7494, 270.7537, 270.7519, 270.7526, 270.7508, 270.7548, 
    270.7515, 270.7556, 270.7552, 270.7541, 270.7518, 270.7513, 270.7507, 
    270.751, 270.7527, 270.753, 270.7541, 270.7545, 270.7553, 270.7561, 
    270.7554, 270.7547, 270.7527, 270.7509, 270.7489, 270.7484, 270.7462, 
    270.748, 270.7451, 270.7477, 270.7431, 270.7512, 270.7477, 270.754, 
    270.7534, 270.7521, 270.7493, 270.7508, 270.749, 270.753, 270.7551, 
    270.7556, 270.7566, 270.7556, 270.7556, 270.7547, 270.755, 270.7526, 
    270.7539, 270.7503, 270.749, 270.7453, 270.743, 270.7407, 270.7397, 
    270.7393, 270.7392 ;

 TREFMXAV_R =
  270.7643, 270.7622, 270.7626, 270.7609, 270.7618, 270.7607, 270.7638, 
    270.7621, 270.7632, 270.7641, 270.7577, 270.7608, 270.7543, 270.7563, 
    270.7512, 270.7546, 270.7505, 270.7512, 270.7488, 270.7495, 270.7466, 
    270.7485, 270.745, 270.747, 270.7467, 270.7486, 270.7601, 270.7581, 
    270.7603, 270.76, 270.7601, 270.7618, 270.7627, 270.7644, 270.7641, 
    270.7628, 270.7598, 270.7608, 270.7583, 270.7583, 270.7555, 270.7568, 
    270.752, 270.7534, 270.7495, 270.7505, 270.7495, 270.7498, 270.7495, 
    270.751, 270.7504, 270.7516, 270.7566, 270.7551, 270.7594, 270.7621, 
    270.7638, 270.765, 270.7648, 270.7645, 270.7628, 270.7612, 270.7599, 
    270.7592, 270.7583, 270.756, 270.7547, 270.7518, 270.7523, 270.7514, 
    270.7506, 270.7492, 270.7494, 270.7488, 270.7514, 270.7497, 270.7526, 
    270.7518, 270.7583, 270.7606, 270.7617, 270.7625, 270.7647, 270.7632, 
    270.7638, 270.7623, 270.7614, 270.7619, 270.7591, 270.7602, 270.7546, 
    270.757, 270.7507, 270.7522, 270.7503, 270.7513, 270.7496, 270.7511, 
    270.7485, 270.748, 270.7484, 270.7469, 270.7512, 270.7495, 270.7619, 
    270.7618, 270.7615, 270.763, 270.7631, 270.7644, 270.7632, 270.7627, 
    270.7614, 270.7606, 270.7599, 270.7582, 270.7565, 270.7539, 270.7521, 
    270.7509, 270.7516, 270.7509, 270.7517, 270.752, 270.7482, 270.7504, 
    270.7471, 270.7473, 270.7488, 270.7473, 270.7618, 270.7622, 270.7636, 
    270.7625, 270.7646, 270.7634, 270.7628, 270.7602, 270.7596, 270.7591, 
    270.7581, 270.7567, 270.7544, 270.7524, 270.7505, 270.7506, 270.7506, 
    270.7502, 270.7512, 270.75, 270.7498, 270.7504, 270.7473, 270.7482, 
    270.7473, 270.7479, 270.7621, 270.7614, 270.7617, 270.761, 270.7615, 
    270.7593, 270.7586, 270.7555, 270.7568, 270.7547, 270.7565, 270.7562, 
    270.7547, 270.7564, 270.7525, 270.7552, 270.7502, 270.7529, 270.75, 
    270.7505, 270.7497, 270.7489, 270.748, 270.7462, 270.7466, 270.7451, 
    270.7603, 270.7594, 270.7595, 270.7585, 270.7578, 270.7563, 270.7538, 
    270.7547, 270.7531, 270.7527, 270.7553, 270.7537, 270.7588, 270.758, 
    270.7585, 270.7602, 270.7546, 270.7575, 270.7521, 270.7536, 270.749, 
    270.7513, 270.7468, 270.7449, 270.7431, 270.741, 270.7589, 270.7595, 
    270.7584, 270.7569, 270.7554, 270.7535, 270.7533, 270.753, 270.7521, 
    270.7513, 270.7529, 270.7511, 270.7579, 270.7543, 270.7597, 270.7581, 
    270.757, 270.7574, 270.7548, 270.7542, 270.7518, 270.753, 270.7454, 
    270.7488, 270.7394, 270.742, 270.7597, 270.7589, 270.756, 270.7574, 
    270.7534, 270.7524, 270.7516, 270.7506, 270.7505, 270.7499, 270.7509, 
    270.75, 270.7535, 270.752, 270.7563, 270.7552, 270.7557, 270.7563, 
    270.7546, 270.7529, 270.7528, 270.7523, 270.7508, 270.7534, 270.7451, 
    270.7503, 270.758, 270.7564, 270.7561, 270.7567, 270.7525, 270.7541, 
    270.7499, 270.7511, 270.7492, 270.7502, 270.7503, 270.7514, 270.7522, 
    270.754, 270.7555, 270.7567, 270.7564, 270.7551, 270.7528, 270.7505, 
    270.751, 270.7494, 270.7537, 270.7519, 270.7526, 270.7508, 270.7548, 
    270.7515, 270.7556, 270.7552, 270.7541, 270.7518, 270.7513, 270.7507, 
    270.751, 270.7527, 270.753, 270.7541, 270.7545, 270.7553, 270.7561, 
    270.7554, 270.7547, 270.7527, 270.7509, 270.7489, 270.7484, 270.7462, 
    270.748, 270.7451, 270.7477, 270.7431, 270.7512, 270.7477, 270.754, 
    270.7534, 270.7521, 270.7493, 270.7508, 270.749, 270.753, 270.7551, 
    270.7556, 270.7566, 270.7556, 270.7556, 270.7547, 270.755, 270.7526, 
    270.7539, 270.7503, 270.749, 270.7453, 270.743, 270.7407, 270.7397, 
    270.7393, 270.7392 ;

 TREFMXAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSA =
  255.2032, 255.203, 255.2031, 255.203, 255.203, 255.2029, 255.2032, 255.203, 
    255.2031, 255.2032, 255.2027, 255.2029, 255.2025, 255.2026, 255.2022, 
    255.2025, 255.2022, 255.2022, 255.2021, 255.2021, 255.2019, 255.202, 
    255.2018, 255.2019, 255.2019, 255.202, 255.2029, 255.2028, 255.2029, 
    255.2029, 255.2029, 255.203, 255.2031, 255.2032, 255.2032, 255.2031, 
    255.2029, 255.2029, 255.2028, 255.2028, 255.2026, 255.2027, 255.2023, 
    255.2024, 255.2021, 255.2022, 255.2021, 255.2021, 255.2021, 255.2022, 
    255.2022, 255.2023, 255.2026, 255.2025, 255.2029, 255.203, 255.2032, 
    255.2032, 255.2032, 255.2032, 255.2031, 255.203, 255.2029, 255.2028, 
    255.2028, 255.2026, 255.2025, 255.2023, 255.2023, 255.2023, 255.2022, 
    255.2021, 255.2021, 255.2021, 255.2023, 255.2021, 255.2023, 255.2023, 
    255.2028, 255.2029, 255.203, 255.2031, 255.2032, 255.2031, 255.2032, 
    255.2031, 255.203, 255.203, 255.2028, 255.2029, 255.2025, 255.2027, 
    255.2022, 255.2023, 255.2022, 255.2022, 255.2021, 255.2022, 255.202, 
    255.202, 255.202, 255.2019, 255.2022, 255.2021, 255.203, 255.203, 
    255.203, 255.2031, 255.2031, 255.2032, 255.2031, 255.2031, 255.203, 
    255.2029, 255.2029, 255.2028, 255.2026, 255.2024, 255.2023, 255.2022, 
    255.2023, 255.2022, 255.2023, 255.2023, 255.202, 255.2022, 255.2019, 
    255.2019, 255.2021, 255.2019, 255.203, 255.203, 255.2032, 255.2031, 
    255.2032, 255.2031, 255.2031, 255.2029, 255.2029, 255.2028, 255.2027, 
    255.2027, 255.2025, 255.2023, 255.2022, 255.2022, 255.2022, 255.2022, 
    255.2022, 255.2021, 255.2021, 255.2022, 255.2019, 255.202, 255.2019, 
    255.202, 255.203, 255.203, 255.203, 255.203, 255.203, 255.2028, 255.2028, 
    255.2026, 255.2027, 255.2025, 255.2026, 255.2026, 255.2025, 255.2026, 
    255.2023, 255.2025, 255.2022, 255.2024, 255.2021, 255.2022, 255.2021, 
    255.2021, 255.202, 255.2019, 255.2019, 255.2018, 255.2029, 255.2029, 
    255.2029, 255.2028, 255.2027, 255.2026, 255.2024, 255.2025, 255.2024, 
    255.2023, 255.2025, 255.2024, 255.2028, 255.2027, 255.2028, 255.2029, 
    255.2025, 255.2027, 255.2023, 255.2024, 255.2021, 255.2022, 255.2019, 
    255.2018, 255.2016, 255.2015, 255.2028, 255.2029, 255.2028, 255.2027, 
    255.2026, 255.2024, 255.2024, 255.2024, 255.2023, 255.2022, 255.2024, 
    255.2022, 255.2027, 255.2025, 255.2029, 255.2028, 255.2027, 255.2027, 
    255.2025, 255.2025, 255.2023, 255.2024, 255.2018, 255.2021, 255.2013, 
    255.2015, 255.2029, 255.2028, 255.2026, 255.2027, 255.2024, 255.2023, 
    255.2023, 255.2022, 255.2022, 255.2021, 255.2022, 255.2021, 255.2024, 
    255.2023, 255.2026, 255.2025, 255.2026, 255.2026, 255.2025, 255.2024, 
    255.2024, 255.2023, 255.2022, 255.2024, 255.2018, 255.2022, 255.2027, 
    255.2026, 255.2026, 255.2027, 255.2023, 255.2025, 255.2021, 255.2022, 
    255.2021, 255.2021, 255.2022, 255.2023, 255.2023, 255.2025, 255.2026, 
    255.2027, 255.2026, 255.2025, 255.2024, 255.2022, 255.2022, 255.2021, 
    255.2024, 255.2023, 255.2023, 255.2022, 255.2025, 255.2023, 255.2026, 
    255.2025, 255.2025, 255.2023, 255.2022, 255.2022, 255.2022, 255.2023, 
    255.2024, 255.2025, 255.2025, 255.2025, 255.2026, 255.2025, 255.2025, 
    255.2023, 255.2022, 255.2021, 255.202, 255.2019, 255.202, 255.2018, 
    255.202, 255.2016, 255.2022, 255.202, 255.2025, 255.2024, 255.2023, 
    255.2021, 255.2022, 255.2021, 255.2024, 255.2025, 255.2026, 255.2026, 
    255.2026, 255.2026, 255.2025, 255.2025, 255.2023, 255.2024, 255.2022, 
    255.2021, 255.2018, 255.2016, 255.2014, 255.2014, 255.2013, 255.2013 ;

 TSAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 TSA_R =
  255.2032, 255.203, 255.2031, 255.203, 255.203, 255.2029, 255.2032, 255.203, 
    255.2031, 255.2032, 255.2027, 255.2029, 255.2025, 255.2026, 255.2022, 
    255.2025, 255.2022, 255.2022, 255.2021, 255.2021, 255.2019, 255.202, 
    255.2018, 255.2019, 255.2019, 255.202, 255.2029, 255.2028, 255.2029, 
    255.2029, 255.2029, 255.203, 255.2031, 255.2032, 255.2032, 255.2031, 
    255.2029, 255.2029, 255.2028, 255.2028, 255.2026, 255.2027, 255.2023, 
    255.2024, 255.2021, 255.2022, 255.2021, 255.2021, 255.2021, 255.2022, 
    255.2022, 255.2023, 255.2026, 255.2025, 255.2029, 255.203, 255.2032, 
    255.2032, 255.2032, 255.2032, 255.2031, 255.203, 255.2029, 255.2028, 
    255.2028, 255.2026, 255.2025, 255.2023, 255.2023, 255.2023, 255.2022, 
    255.2021, 255.2021, 255.2021, 255.2023, 255.2021, 255.2023, 255.2023, 
    255.2028, 255.2029, 255.203, 255.2031, 255.2032, 255.2031, 255.2032, 
    255.2031, 255.203, 255.203, 255.2028, 255.2029, 255.2025, 255.2027, 
    255.2022, 255.2023, 255.2022, 255.2022, 255.2021, 255.2022, 255.202, 
    255.202, 255.202, 255.2019, 255.2022, 255.2021, 255.203, 255.203, 
    255.203, 255.2031, 255.2031, 255.2032, 255.2031, 255.2031, 255.203, 
    255.2029, 255.2029, 255.2028, 255.2026, 255.2024, 255.2023, 255.2022, 
    255.2023, 255.2022, 255.2023, 255.2023, 255.202, 255.2022, 255.2019, 
    255.2019, 255.2021, 255.2019, 255.203, 255.203, 255.2032, 255.2031, 
    255.2032, 255.2031, 255.2031, 255.2029, 255.2029, 255.2028, 255.2027, 
    255.2027, 255.2025, 255.2023, 255.2022, 255.2022, 255.2022, 255.2022, 
    255.2022, 255.2021, 255.2021, 255.2022, 255.2019, 255.202, 255.2019, 
    255.202, 255.203, 255.203, 255.203, 255.203, 255.203, 255.2028, 255.2028, 
    255.2026, 255.2027, 255.2025, 255.2026, 255.2026, 255.2025, 255.2026, 
    255.2023, 255.2025, 255.2022, 255.2024, 255.2021, 255.2022, 255.2021, 
    255.2021, 255.202, 255.2019, 255.2019, 255.2018, 255.2029, 255.2029, 
    255.2029, 255.2028, 255.2027, 255.2026, 255.2024, 255.2025, 255.2024, 
    255.2023, 255.2025, 255.2024, 255.2028, 255.2027, 255.2028, 255.2029, 
    255.2025, 255.2027, 255.2023, 255.2024, 255.2021, 255.2022, 255.2019, 
    255.2018, 255.2016, 255.2015, 255.2028, 255.2029, 255.2028, 255.2027, 
    255.2026, 255.2024, 255.2024, 255.2024, 255.2023, 255.2022, 255.2024, 
    255.2022, 255.2027, 255.2025, 255.2029, 255.2028, 255.2027, 255.2027, 
    255.2025, 255.2025, 255.2023, 255.2024, 255.2018, 255.2021, 255.2013, 
    255.2015, 255.2029, 255.2028, 255.2026, 255.2027, 255.2024, 255.2023, 
    255.2023, 255.2022, 255.2022, 255.2021, 255.2022, 255.2021, 255.2024, 
    255.2023, 255.2026, 255.2025, 255.2026, 255.2026, 255.2025, 255.2024, 
    255.2024, 255.2023, 255.2022, 255.2024, 255.2018, 255.2022, 255.2027, 
    255.2026, 255.2026, 255.2027, 255.2023, 255.2025, 255.2021, 255.2022, 
    255.2021, 255.2021, 255.2022, 255.2023, 255.2023, 255.2025, 255.2026, 
    255.2027, 255.2026, 255.2025, 255.2024, 255.2022, 255.2022, 255.2021, 
    255.2024, 255.2023, 255.2023, 255.2022, 255.2025, 255.2023, 255.2026, 
    255.2025, 255.2025, 255.2023, 255.2022, 255.2022, 255.2022, 255.2023, 
    255.2024, 255.2025, 255.2025, 255.2025, 255.2026, 255.2025, 255.2025, 
    255.2023, 255.2022, 255.2021, 255.202, 255.2019, 255.202, 255.2018, 
    255.202, 255.2016, 255.2022, 255.202, 255.2025, 255.2024, 255.2023, 
    255.2021, 255.2022, 255.2021, 255.2024, 255.2025, 255.2026, 255.2026, 
    255.2026, 255.2026, 255.2025, 255.2025, 255.2023, 255.2024, 255.2022, 
    255.2021, 255.2018, 255.2016, 255.2014, 255.2014, 255.2013, 255.2013 ;

 TSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSOI =
  253.6898, 253.6917, 253.6913, 253.6929, 253.692, 253.693, 253.6902, 
    253.6918, 253.6908, 253.69, 253.6958, 253.6929, 253.6988, 253.697, 
    253.7016, 253.6985, 253.7023, 253.7016, 253.7037, 253.7031, 253.7058, 
    253.704, 253.7072, 253.7054, 253.7057, 253.7039, 253.6935, 253.6954, 
    253.6934, 253.6937, 253.6936, 253.692, 253.6913, 253.6897, 253.69, 
    253.6911, 253.6938, 253.6929, 253.6952, 253.6952, 253.6977, 253.6966, 
    253.7008, 253.6996, 253.7031, 253.7023, 253.7031, 253.7028, 253.7031, 
    253.7018, 253.7023, 253.7012, 253.6968, 253.6981, 253.6942, 253.6918, 
    253.6903, 253.6892, 253.6893, 253.6896, 253.6911, 253.6926, 253.6937, 
    253.6944, 253.6952, 253.6973, 253.6985, 253.701, 253.7006, 253.7014, 
    253.7022, 253.7034, 253.7032, 253.7038, 253.7014, 253.703, 253.7004, 
    253.7011, 253.6952, 253.6932, 253.6922, 253.6914, 253.6895, 253.6908, 
    253.6903, 253.6916, 253.6924, 253.692, 253.6945, 253.6935, 253.6985, 
    253.6964, 253.7021, 253.7007, 253.7024, 253.7015, 253.703, 253.7017, 
    253.704, 253.7045, 253.7041, 253.7055, 253.7016, 253.7031, 253.692, 
    253.692, 253.6923, 253.691, 253.6909, 253.6897, 253.6908, 253.6912, 
    253.6924, 253.6931, 253.6938, 253.6953, 253.6969, 253.6991, 253.7008, 
    253.7019, 253.7012, 253.7018, 253.7012, 253.7009, 253.7043, 253.7023, 
    253.7053, 253.7051, 253.7038, 253.7051, 253.6921, 253.6917, 253.6904, 
    253.6914, 253.6895, 253.6906, 253.6912, 253.6935, 253.694, 253.6945, 
    253.6954, 253.6966, 253.6987, 253.7005, 253.7022, 253.7021, 253.7021, 
    253.7025, 253.7016, 253.7027, 253.7028, 253.7024, 253.7051, 253.7043, 
    253.7051, 253.7046, 253.6918, 253.6925, 253.6921, 253.6927, 253.6923, 
    253.6943, 253.6949, 253.6977, 253.6966, 253.6984, 253.6968, 253.6971, 
    253.6984, 253.6969, 253.7004, 253.698, 253.7025, 253.7, 253.7027, 
    253.7022, 253.703, 253.7037, 253.7045, 253.7061, 253.7058, 253.7071, 
    253.6934, 253.6942, 253.6942, 253.695, 253.6956, 253.697, 253.6992, 
    253.6984, 253.6999, 253.7002, 253.6979, 253.6993, 253.6948, 253.6955, 
    253.6951, 253.6935, 253.6986, 253.6959, 253.7008, 253.6994, 253.7036, 
    253.7015, 253.7056, 253.7072, 253.709, 253.7108, 253.6947, 253.6941, 
    253.6951, 253.6965, 253.6978, 253.6995, 253.6997, 253.7, 253.7008, 
    253.7015, 253.7001, 253.7017, 253.6956, 253.6988, 253.6939, 253.6953, 
    253.6964, 253.696, 253.6983, 253.6989, 253.7011, 253.7, 253.7068, 
    253.7038, 253.7123, 253.7099, 253.6939, 253.6947, 253.6973, 253.696, 
    253.6996, 253.7005, 253.7012, 253.7021, 253.7022, 253.7027, 253.7019, 
    253.7027, 253.6995, 253.7009, 253.697, 253.6979, 253.6975, 253.697, 
    253.6985, 253.7001, 253.7001, 253.7006, 253.702, 253.6996, 253.7071, 
    253.7024, 253.6955, 253.6969, 253.6971, 253.6966, 253.7004, 253.699, 
    253.7027, 253.7017, 253.7034, 253.7025, 253.7024, 253.7014, 253.7007, 
    253.6991, 253.6977, 253.6967, 253.6969, 253.6981, 253.7002, 253.7022, 
    253.7018, 253.7032, 253.6994, 253.701, 253.7003, 253.702, 253.6984, 
    253.7013, 253.6976, 253.698, 253.699, 253.701, 253.7016, 253.702, 
    253.7018, 253.7002, 253.7, 253.699, 253.6987, 253.6979, 253.6972, 
    253.6978, 253.6984, 253.7003, 253.7019, 253.7037, 253.7041, 253.7061, 
    253.7044, 253.7072, 253.7048, 253.7089, 253.7016, 253.7048, 253.699, 
    253.6997, 253.7008, 253.7033, 253.702, 253.7036, 253.7, 253.6981, 
    253.6976, 253.6967, 253.6977, 253.6976, 253.6985, 253.6982, 253.7003, 
    253.6992, 253.7024, 253.7036, 253.707, 253.709, 253.7111, 253.7121, 
    253.7124, 253.7125,
  255.2211, 255.2229, 255.2225, 255.2239, 255.2232, 255.2241, 255.2215, 
    255.2229, 255.222, 255.2213, 255.2266, 255.224, 255.2295, 255.2278, 
    255.2321, 255.2292, 255.2327, 255.232, 255.2341, 255.2335, 255.236, 
    255.2343, 255.2374, 255.2356, 255.2359, 255.2343, 255.2245, 255.2263, 
    255.2244, 255.2247, 255.2246, 255.2232, 255.2224, 255.221, 255.2212, 
    255.2223, 255.2248, 255.224, 255.2261, 255.2261, 255.2284, 255.2274, 
    255.2313, 255.2302, 255.2335, 255.2327, 255.2335, 255.2332, 255.2335, 
    255.2322, 255.2328, 255.2317, 255.2276, 255.2288, 255.2251, 255.2229, 
    255.2215, 255.2205, 255.2206, 255.2209, 255.2223, 255.2237, 255.2247, 
    255.2254, 255.2261, 255.228, 255.2291, 255.2316, 255.2311, 255.2319, 
    255.2326, 255.2338, 255.2336, 255.2341, 255.2319, 255.2333, 255.2309, 
    255.2316, 255.2261, 255.2242, 255.2233, 255.2226, 255.2207, 255.222, 
    255.2215, 255.2227, 255.2235, 255.2231, 255.2254, 255.2245, 255.2292, 
    255.2272, 255.2325, 255.2312, 255.2328, 255.232, 255.2334, 255.2321, 
    255.2343, 255.2348, 255.2345, 255.2357, 255.2321, 255.2334, 255.2231, 
    255.2231, 255.2234, 255.2222, 255.2221, 255.221, 255.222, 255.2224, 
    255.2235, 255.2242, 255.2248, 255.2261, 255.2276, 255.2298, 255.2313, 
    255.2323, 255.2317, 255.2323, 255.2316, 255.2314, 255.2346, 255.2328, 
    255.2355, 255.2354, 255.2341, 255.2354, 255.2232, 255.2228, 255.2216, 
    255.2226, 255.2208, 255.2218, 255.2223, 255.2245, 255.225, 255.2254, 
    255.2263, 255.2274, 255.2294, 255.231, 255.2326, 255.2325, 255.2326, 
    255.2329, 255.232, 255.233, 255.2332, 255.2328, 255.2354, 255.2346, 
    255.2354, 255.2349, 255.2229, 255.2235, 255.2232, 255.2238, 255.2234, 
    255.2252, 255.2258, 255.2284, 255.2274, 255.2291, 255.2276, 255.2278, 
    255.2291, 255.2276, 255.2309, 255.2287, 255.2329, 255.2306, 255.2331, 
    255.2326, 255.2334, 255.234, 255.2348, 255.2363, 255.236, 255.2372, 
    255.2244, 255.2252, 255.2251, 255.2259, 255.2265, 255.2278, 255.2298, 
    255.2291, 255.2305, 255.2308, 255.2286, 255.2299, 255.2257, 255.2263, 
    255.226, 255.2245, 255.2292, 255.2268, 255.2313, 255.23, 255.2339, 
    255.2319, 255.2358, 255.2374, 255.239, 255.2407, 255.2256, 255.2251, 
    255.226, 255.2273, 255.2285, 255.2301, 255.2303, 255.2305, 255.2313, 
    255.232, 255.2306, 255.2321, 255.2265, 255.2294, 255.2249, 255.2262, 
    255.2272, 255.2268, 255.229, 255.2295, 255.2316, 255.2305, 255.237, 
    255.2341, 255.2421, 255.2399, 255.2249, 255.2256, 255.228, 255.2269, 
    255.2302, 255.231, 255.2317, 255.2325, 255.2326, 255.2331, 255.2323, 
    255.2331, 255.2301, 255.2314, 255.2278, 255.2286, 255.2282, 255.2278, 
    255.2292, 255.2306, 255.2307, 255.2312, 255.2324, 255.2302, 255.2373, 
    255.2328, 255.2264, 255.2277, 255.2279, 255.2274, 255.2309, 255.2296, 
    255.2331, 255.2322, 255.2337, 255.233, 255.2328, 255.2319, 255.2312, 
    255.2297, 255.2284, 255.2275, 255.2277, 255.2288, 255.2307, 255.2326, 
    255.2322, 255.2336, 255.2299, 255.2315, 255.2309, 255.2324, 255.229, 
    255.2318, 255.2283, 255.2286, 255.2296, 255.2315, 255.232, 255.2325, 
    255.2322, 255.2308, 255.2306, 255.2296, 255.2293, 255.2286, 255.228, 
    255.2285, 255.2291, 255.2308, 255.2323, 255.234, 255.2344, 255.2363, 
    255.2347, 255.2373, 255.235, 255.239, 255.232, 255.235, 255.2297, 
    255.2303, 255.2313, 255.2337, 255.2324, 255.2339, 255.2306, 255.2288, 
    255.2284, 255.2275, 255.2284, 255.2283, 255.2291, 255.2289, 255.2309, 
    255.2298, 255.2328, 255.2339, 255.2371, 255.239, 255.241, 255.2419, 
    255.2422, 255.2423,
  257.287, 257.2885, 257.2882, 257.2893, 257.2887, 257.2894, 257.2874, 
    257.2885, 257.2878, 257.2872, 257.2915, 257.2894, 257.2938, 257.2924, 
    257.2959, 257.2936, 257.2964, 257.2959, 257.2975, 257.2971, 257.2991, 
    257.2978, 257.3003, 257.2988, 257.299, 257.2977, 257.2898, 257.2912, 
    257.2897, 257.2899, 257.2899, 257.2887, 257.2881, 257.287, 257.2872, 
    257.288, 257.29, 257.2894, 257.2911, 257.291, 257.293, 257.2921, 
    257.2953, 257.2944, 257.2971, 257.2964, 257.2971, 257.2969, 257.2971, 
    257.2961, 257.2965, 257.2956, 257.2922, 257.2932, 257.2903, 257.2885, 
    257.2874, 257.2866, 257.2867, 257.2869, 257.288, 257.2891, 257.2899, 
    257.2905, 257.291, 257.2926, 257.2935, 257.2955, 257.2952, 257.2957, 
    257.2964, 257.2973, 257.2971, 257.2976, 257.2957, 257.297, 257.295, 
    257.2955, 257.2911, 257.2896, 257.2888, 257.2882, 257.2868, 257.2878, 
    257.2874, 257.2884, 257.2889, 257.2887, 257.2905, 257.2898, 257.2936, 
    257.2919, 257.2963, 257.2952, 257.2965, 257.2959, 257.297, 257.296, 
    257.2978, 257.2981, 257.2979, 257.2989, 257.2959, 257.2971, 257.2886, 
    257.2887, 257.2889, 257.2879, 257.2878, 257.287, 257.2878, 257.2881, 
    257.289, 257.2895, 257.29, 257.2911, 257.2923, 257.294, 257.2953, 
    257.2961, 257.2956, 257.2961, 257.2956, 257.2953, 257.298, 257.2965, 
    257.2987, 257.2986, 257.2976, 257.2986, 257.2887, 257.2885, 257.2875, 
    257.2882, 257.2869, 257.2876, 257.2881, 257.2898, 257.2902, 257.2905, 
    257.2912, 257.2921, 257.2937, 257.2951, 257.2964, 257.2963, 257.2963, 
    257.2966, 257.2959, 257.2967, 257.2968, 257.2965, 257.2986, 257.298, 
    257.2986, 257.2982, 257.2885, 257.289, 257.2888, 257.2892, 257.2889, 
    257.2904, 257.2908, 257.293, 257.2921, 257.2935, 257.2923, 257.2925, 
    257.2935, 257.2923, 257.295, 257.2932, 257.2966, 257.2947, 257.2967, 
    257.2964, 257.297, 257.2975, 257.2982, 257.2994, 257.2991, 257.3001, 
    257.2897, 257.2903, 257.2903, 257.2909, 257.2914, 257.2924, 257.2941, 
    257.2935, 257.2946, 257.2949, 257.2931, 257.2942, 257.2907, 257.2913, 
    257.291, 257.2898, 257.2936, 257.2916, 257.2953, 257.2943, 257.2974, 
    257.2958, 257.299, 257.3003, 257.3016, 257.303, 257.2907, 257.2903, 
    257.291, 257.292, 257.293, 257.2943, 257.2944, 257.2947, 257.2953, 
    257.2958, 257.2947, 257.296, 257.2914, 257.2938, 257.2901, 257.2912, 
    257.292, 257.2916, 257.2934, 257.2939, 257.2955, 257.2947, 257.2999, 
    257.2976, 257.3042, 257.3023, 257.2901, 257.2907, 257.2926, 257.2917, 
    257.2944, 257.295, 257.2956, 257.2963, 257.2964, 257.2968, 257.2961, 
    257.2968, 257.2943, 257.2954, 257.2924, 257.2931, 257.2928, 257.2924, 
    257.2936, 257.2948, 257.2948, 257.2952, 257.2962, 257.2944, 257.3002, 
    257.2966, 257.2913, 257.2924, 257.2925, 257.2921, 257.295, 257.2939, 
    257.2968, 257.296, 257.2973, 257.2966, 257.2965, 257.2957, 257.2953, 
    257.294, 257.293, 257.2922, 257.2924, 257.2932, 257.2948, 257.2964, 
    257.296, 257.2972, 257.2942, 257.2954, 257.295, 257.2962, 257.2935, 
    257.2957, 257.2929, 257.2932, 257.2939, 257.2955, 257.2959, 257.2963, 
    257.296, 257.2949, 257.2947, 257.2939, 257.2937, 257.2931, 257.2926, 
    257.293, 257.2935, 257.2949, 257.2961, 257.2975, 257.2979, 257.2994, 
    257.2981, 257.3002, 257.2984, 257.3016, 257.2959, 257.2983, 257.294, 
    257.2944, 257.2953, 257.2972, 257.2962, 257.2975, 257.2947, 257.2932, 
    257.2929, 257.2922, 257.2929, 257.2929, 257.2935, 257.2933, 257.295, 
    257.2941, 257.2965, 257.2975, 257.3, 257.3016, 257.3033, 257.304, 
    257.3042, 257.3043,
  259.794, 259.7949, 259.7947, 259.7953, 259.795, 259.7954, 259.7942, 
    259.7949, 259.7944, 259.7941, 259.7966, 259.7954, 259.798, 259.7972, 
    259.7993, 259.7979, 259.7996, 259.7993, 259.8002, 259.8, 259.8012, 
    259.8004, 259.8019, 259.801, 259.8011, 259.8004, 259.7957, 259.7965, 
    259.7956, 259.7957, 259.7957, 259.795, 259.7946, 259.794, 259.7941, 
    259.7946, 259.7958, 259.7954, 259.7964, 259.7964, 259.7975, 259.797, 
    259.7989, 259.7984, 259.8, 259.7996, 259.8, 259.7998, 259.8, 259.7993, 
    259.7996, 259.7991, 259.7971, 259.7976, 259.7959, 259.7949, 259.7942, 
    259.7938, 259.7938, 259.7939, 259.7946, 259.7952, 259.7957, 259.7961, 
    259.7964, 259.7973, 259.7978, 259.799, 259.7988, 259.7992, 259.7995, 
    259.8001, 259.8, 259.8003, 259.7992, 259.7999, 259.7987, 259.799, 
    259.7964, 259.7955, 259.795, 259.7947, 259.7939, 259.7945, 259.7942, 
    259.7948, 259.7951, 259.795, 259.7961, 259.7956, 259.7979, 259.7969, 
    259.7995, 259.7989, 259.7996, 259.7992, 259.7999, 259.7993, 259.8004, 
    259.8006, 259.8004, 259.8011, 259.7993, 259.7999, 259.795, 259.795, 
    259.7951, 259.7945, 259.7945, 259.794, 259.7944, 259.7946, 259.7952, 
    259.7955, 259.7957, 259.7964, 259.7971, 259.7981, 259.7989, 259.7994, 
    259.7991, 259.7993, 259.799, 259.7989, 259.8005, 259.7996, 259.801, 
    259.8009, 259.8003, 259.8009, 259.795, 259.7948, 259.7943, 259.7947, 
    259.7939, 259.7943, 259.7946, 259.7956, 259.7959, 259.7961, 259.7965, 
    259.797, 259.7979, 259.7988, 259.7995, 259.7995, 259.7995, 259.7997, 
    259.7993, 259.7997, 259.7998, 259.7996, 259.8009, 259.8005, 259.8009, 
    259.8007, 259.7949, 259.7952, 259.795, 259.7953, 259.7951, 259.796, 
    259.7962, 259.7975, 259.797, 259.7978, 259.7971, 259.7972, 259.7978, 
    259.7971, 259.7987, 259.7976, 259.7997, 259.7986, 259.7997, 259.7995, 
    259.7999, 259.8002, 259.8006, 259.8014, 259.8012, 259.8018, 259.7956, 
    259.7959, 259.7959, 259.7963, 259.7966, 259.7972, 259.7982, 259.7978, 
    259.7985, 259.7986, 259.7976, 259.7982, 259.7962, 259.7965, 259.7963, 
    259.7956, 259.7979, 259.7967, 259.7989, 259.7982, 259.8002, 259.7992, 
    259.8011, 259.8019, 259.8027, 259.8036, 259.7961, 259.7959, 259.7964, 
    259.7969, 259.7975, 259.7983, 259.7984, 259.7985, 259.7989, 259.7992, 
    259.7986, 259.7993, 259.7966, 259.798, 259.7958, 259.7964, 259.7969, 
    259.7967, 259.7978, 259.798, 259.799, 259.7985, 259.8017, 259.8003, 
    259.8043, 259.8032, 259.7958, 259.7961, 259.7973, 259.7968, 259.7983, 
    259.7987, 259.7991, 259.7995, 259.7995, 259.7998, 259.7994, 259.7998, 
    259.7983, 259.799, 259.7972, 259.7976, 259.7974, 259.7972, 259.7979, 
    259.7986, 259.7986, 259.7988, 259.7994, 259.7984, 259.8018, 259.7997, 
    259.7965, 259.7971, 259.7972, 259.797, 259.7987, 259.7981, 259.7998, 
    259.7993, 259.8001, 259.7997, 259.7997, 259.7992, 259.7989, 259.7981, 
    259.7975, 259.797, 259.7971, 259.7977, 259.7986, 259.7995, 259.7993, 
    259.8, 259.7982, 259.799, 259.7987, 259.7994, 259.7978, 259.7992, 
    259.7975, 259.7976, 259.7981, 259.799, 259.7992, 259.7995, 259.7993, 
    259.7986, 259.7985, 259.7981, 259.7979, 259.7976, 259.7973, 259.7975, 
    259.7978, 259.7986, 259.7994, 259.8002, 259.8004, 259.8014, 259.8006, 
    259.8018, 259.8007, 259.8027, 259.7993, 259.8007, 259.7981, 259.7984, 
    259.7989, 259.8001, 259.7994, 259.8002, 259.7985, 259.7977, 259.7975, 
    259.7971, 259.7975, 259.7975, 259.7979, 259.7977, 259.7987, 259.7982, 
    259.7996, 259.8002, 259.8018, 259.8027, 259.8037, 259.8042, 259.8043, 
    259.8044,
  262.0097, 262.0099, 262.0099, 262.0101, 262.01, 262.0101, 262.0098, 
    262.0099, 262.0098, 262.0097, 262.0104, 262.0101, 262.0108, 262.0106, 
    262.0111, 262.0107, 262.0112, 262.0111, 262.0114, 262.0113, 262.0117, 
    262.0114, 262.0119, 262.0116, 262.0117, 262.0114, 262.0101, 262.0103, 
    262.0101, 262.0102, 262.0101, 262.01, 262.0099, 262.0097, 262.0097, 
    262.0099, 262.0102, 262.0101, 262.0103, 262.0103, 262.0106, 262.0105, 
    262.011, 262.0109, 262.0113, 262.0112, 262.0113, 262.0113, 262.0113, 
    262.0111, 262.0112, 262.0111, 262.0105, 262.0107, 262.0102, 262.0099, 
    262.0098, 262.0096, 262.0097, 262.0097, 262.0099, 262.01, 262.0102, 
    262.0103, 262.0103, 262.0106, 262.0107, 262.011, 262.011, 262.0111, 
    262.0112, 262.0114, 262.0113, 262.0114, 262.0111, 262.0113, 262.011, 
    262.011, 262.0103, 262.0101, 262.01, 262.0099, 262.0097, 262.0098, 
    262.0098, 262.0099, 262.01, 262.0099, 262.0103, 262.0101, 262.0107, 
    262.0105, 262.0112, 262.011, 262.0112, 262.0111, 262.0113, 262.0111, 
    262.0114, 262.0115, 262.0114, 262.0116, 262.0111, 262.0113, 262.0099, 
    262.01, 262.01, 262.0099, 262.0098, 262.0097, 262.0098, 262.0099, 262.01, 
    262.0101, 262.0102, 262.0103, 262.0105, 262.0108, 262.011, 262.0112, 
    262.0111, 262.0111, 262.0111, 262.011, 262.0115, 262.0112, 262.0116, 
    262.0116, 262.0114, 262.0116, 262.01, 262.0099, 262.0098, 262.0099, 
    262.0097, 262.0098, 262.0099, 262.0101, 262.0102, 262.0103, 262.0103, 
    262.0105, 262.0107, 262.011, 262.0112, 262.0112, 262.0112, 262.0112, 
    262.0111, 262.0113, 262.0113, 262.0112, 262.0116, 262.0115, 262.0116, 
    262.0115, 262.0099, 262.01, 262.01, 262.01, 262.01, 262.0102, 262.0103, 
    262.0106, 262.0105, 262.0107, 262.0105, 262.0106, 262.0107, 262.0105, 
    262.011, 262.0107, 262.0112, 262.0109, 262.0113, 262.0112, 262.0113, 
    262.0114, 262.0115, 262.0117, 262.0117, 262.0119, 262.0101, 262.0102, 
    262.0102, 262.0103, 262.0104, 262.0106, 262.0108, 262.0107, 262.0109, 
    262.011, 262.0107, 262.0108, 262.0103, 262.0104, 262.0103, 262.0101, 
    262.0107, 262.0104, 262.011, 262.0108, 262.0114, 262.0111, 262.0117, 
    262.0119, 262.0121, 262.0124, 262.0103, 262.0102, 262.0103, 262.0105, 
    262.0107, 262.0109, 262.0109, 262.0109, 262.011, 262.0111, 262.0109, 
    262.0111, 262.0104, 262.0108, 262.0102, 262.0103, 262.0105, 262.0104, 
    262.0107, 262.0108, 262.011, 262.0109, 262.0118, 262.0114, 262.0126, 
    262.0123, 262.0102, 262.0103, 262.0106, 262.0104, 262.0109, 262.011, 
    262.0111, 262.0112, 262.0112, 262.0113, 262.0112, 262.0113, 262.0109, 
    262.011, 262.0106, 262.0107, 262.0106, 262.0106, 262.0107, 262.0109, 
    262.0109, 262.011, 262.0112, 262.0109, 262.0119, 262.0112, 262.0104, 
    262.0105, 262.0106, 262.0105, 262.011, 262.0108, 262.0113, 262.0111, 
    262.0114, 262.0112, 262.0112, 262.0111, 262.011, 262.0108, 262.0106, 
    262.0105, 262.0105, 262.0107, 262.0109, 262.0112, 262.0111, 262.0113, 
    262.0108, 262.011, 262.011, 262.0112, 262.0107, 262.0111, 262.0106, 
    262.0107, 262.0108, 262.011, 262.0111, 262.0112, 262.0111, 262.011, 
    262.0109, 262.0108, 262.0107, 262.0107, 262.0106, 262.0107, 262.0107, 
    262.011, 262.0112, 262.0114, 262.0114, 262.0117, 262.0115, 262.0119, 
    262.0115, 262.0121, 262.0111, 262.0115, 262.0108, 262.0109, 262.011, 
    262.0114, 262.0112, 262.0114, 262.0109, 262.0107, 262.0106, 262.0105, 
    262.0106, 262.0106, 262.0107, 262.0107, 262.011, 262.0108, 262.0112, 
    262.0114, 262.0118, 262.0121, 262.0125, 262.0126, 262.0126, 262.0126,
  262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 262.9985, 
    262.9985, 262.9985,
  263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 263.1447, 
    263.1447, 263.1447,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15 ;

 TSOI_10CM =
  263.2749, 263.2867, 263.2844, 263.2939, 263.2887, 263.2949, 263.2773, 
    263.2872, 263.2809, 263.276, 263.3123, 263.2944, 263.3308, 263.3195, 
    263.3478, 263.329, 263.3516, 263.3473, 263.3603, 263.3566, 263.3732, 
    263.362, 263.3818, 263.3705, 263.3723, 263.3617, 263.298, 263.3101, 
    263.2973, 263.299, 263.2982, 263.2888, 263.284, 263.274, 263.2758, 
    263.2832, 263.2998, 263.2942, 263.3083, 263.308, 263.3237, 263.3167, 
    263.3428, 263.3354, 263.3568, 263.3514, 263.3565, 263.3549, 263.3565, 
    263.3486, 263.352, 263.3451, 263.318, 263.326, 263.302, 263.2874, 
    263.2778, 263.2709, 263.2719, 263.2737, 263.2832, 263.2921, 263.299, 
    263.3035, 263.308, 263.3214, 263.3285, 263.3442, 263.3414, 263.3462, 
    263.3508, 263.3586, 263.3573, 263.3607, 263.3461, 263.3558, 263.3398, 
    263.3442, 263.3091, 263.2957, 263.2899, 263.2849, 263.2726, 263.2811, 
    263.2777, 263.2857, 263.2907, 263.2882, 263.3036, 263.2976, 263.3289, 
    263.3156, 263.3503, 263.342, 263.3523, 263.347, 263.356, 263.3479, 
    263.3619, 263.365, 263.3629, 263.3709, 263.3475, 263.3565, 263.2882, 
    263.2886, 263.2905, 263.2821, 263.2816, 263.274, 263.2808, 263.2837, 
    263.291, 263.2954, 263.2995, 263.3086, 263.3186, 263.3326, 263.3425, 
    263.3492, 263.3451, 263.3488, 263.3447, 263.3428, 263.3638, 263.352, 
    263.3698, 263.3688, 263.3607, 263.3689, 263.2888, 263.2865, 263.2784, 
    263.2848, 263.2732, 263.2796, 263.2834, 263.2978, 263.3009, 263.3039, 
    263.3096, 263.317, 263.3299, 263.3409, 263.3511, 263.3504, 263.3506, 
    263.3529, 263.3473, 263.3538, 263.3549, 263.3521, 263.3686, 263.3639, 
    263.3687, 263.3657, 263.2873, 263.2912, 263.2891, 263.2931, 263.2903, 
    263.3028, 263.3065, 263.324, 263.3169, 263.3282, 263.3181, 263.3199, 
    263.3285, 263.3186, 263.3403, 263.3256, 263.353, 263.3383, 263.3539, 
    263.3511, 263.3557, 263.36, 263.3652, 263.3749, 263.3727, 263.3808, 
    263.2971, 263.3022, 263.3018, 263.3071, 263.311, 263.3195, 263.333, 
    263.328, 263.3373, 263.3391, 263.325, 263.3337, 263.3056, 263.3102, 
    263.3075, 263.2975, 263.3291, 263.313, 263.3427, 263.334, 263.3593, 
    263.3467, 263.3715, 263.382, 263.3919, 263.4034, 263.305, 263.3015, 
    263.3077, 263.3163, 263.3242, 263.3346, 263.3356, 263.3376, 263.3426, 
    263.3468, 263.3382, 263.3479, 263.3112, 263.3305, 263.3002, 263.3094, 
    263.3158, 263.313, 263.3274, 263.3308, 263.3444, 263.3374, 263.3794, 
    263.3608, 263.4122, 263.3979, 263.3003, 263.305, 263.3211, 263.3135, 
    263.3353, 263.3406, 263.3449, 263.3504, 263.351, 263.3543, 263.349, 
    263.3541, 263.3346, 263.3433, 263.3193, 263.3252, 263.3225, 263.3195, 
    263.3286, 263.3383, 263.3386, 263.3416, 263.3503, 263.3354, 263.3817, 
    263.3531, 263.3101, 263.319, 263.3203, 263.3168, 263.3401, 263.3317, 
    263.3542, 263.3481, 263.3582, 263.3532, 263.3524, 263.3461, 263.3421, 
    263.3321, 263.3239, 263.3173, 263.3189, 263.326, 263.3389, 263.3511, 
    263.3484, 263.3574, 263.3337, 263.3436, 263.3398, 263.3498, 263.3279, 
    263.3465, 263.3231, 263.3251, 263.3315, 263.3443, 263.3471, 263.3502, 
    263.3483, 263.3392, 263.3378, 263.3314, 263.3296, 263.3247, 263.3206, 
    263.3243, 263.3282, 263.3393, 263.3492, 263.36, 263.3627, 263.3752, 
    263.365, 263.3819, 263.3674, 263.3924, 263.3476, 263.3671, 263.3318, 
    263.3356, 263.3425, 263.3582, 263.3498, 263.3597, 263.3377, 263.3262, 
    263.3233, 263.3177, 263.3234, 263.323, 263.3284, 263.3266, 263.3396, 
    263.3327, 263.3524, 263.3596, 263.38, 263.3924, 263.4051, 263.4106, 
    263.4124, 263.4131 ;

 TSOI_ICE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TV =
  253.9098, 253.9106, 253.9105, 253.9111, 253.9108, 253.9112, 253.91, 
    253.9107, 253.9102, 253.9099, 253.9124, 253.9112, 253.9138, 253.913, 
    253.9151, 253.9137, 253.9153, 253.915, 253.916, 253.9157, 253.9169, 
    253.9161, 253.9175, 253.9167, 253.9168, 253.9161, 253.9115, 253.9123, 
    253.9114, 253.9115, 253.9115, 253.9108, 253.9104, 253.9097, 253.9099, 
    253.9104, 253.9116, 253.9112, 253.9122, 253.9122, 253.9133, 253.9128, 
    253.9147, 253.9142, 253.9157, 253.9153, 253.9157, 253.9156, 253.9157, 
    253.9151, 253.9154, 253.9149, 253.9129, 253.9135, 253.9117, 253.9107, 
    253.91, 253.9095, 253.9096, 253.9097, 253.9104, 253.911, 253.9115, 
    253.9118, 253.9122, 253.9131, 253.9137, 253.9148, 253.9146, 253.9149, 
    253.9153, 253.9158, 253.9158, 253.916, 253.9149, 253.9156, 253.9145, 
    253.9148, 253.9122, 253.9113, 253.9108, 253.9105, 253.9096, 253.9102, 
    253.91, 253.9106, 253.9109, 253.9108, 253.9119, 253.9114, 253.9137, 
    253.9127, 253.9153, 253.9146, 253.9154, 253.915, 253.9157, 253.9151, 
    253.9161, 253.9163, 253.9162, 253.9168, 253.9151, 253.9157, 253.9107, 
    253.9108, 253.9109, 253.9103, 253.9103, 253.9097, 253.9102, 253.9104, 
    253.9109, 253.9113, 253.9116, 253.9122, 253.9129, 253.914, 253.9147, 
    253.9152, 253.9149, 253.9151, 253.9148, 253.9147, 253.9162, 253.9154, 
    253.9167, 253.9166, 253.916, 253.9166, 253.9108, 253.9106, 253.91, 
    253.9105, 253.9097, 253.9101, 253.9104, 253.9114, 253.9117, 253.9119, 
    253.9123, 253.9128, 253.9138, 253.9146, 253.9153, 253.9153, 253.9153, 
    253.9154, 253.915, 253.9155, 253.9156, 253.9154, 253.9166, 253.9162, 
    253.9166, 253.9164, 253.9107, 253.911, 253.9108, 253.9111, 253.9109, 
    253.9118, 253.912, 253.9133, 253.9128, 253.9136, 253.9129, 253.913, 
    253.9136, 253.9129, 253.9145, 253.9134, 253.9155, 253.9144, 253.9155, 
    253.9153, 253.9156, 253.916, 253.9164, 253.9171, 253.9169, 253.9175, 
    253.9114, 253.9117, 253.9117, 253.9121, 253.9124, 253.913, 253.914, 
    253.9136, 253.9143, 253.9144, 253.9134, 253.914, 253.912, 253.9123, 
    253.9121, 253.9114, 253.9137, 253.9125, 253.9147, 253.9141, 253.9159, 
    253.915, 253.9168, 253.9175, 253.9183, 253.9191, 253.912, 253.9117, 
    253.9122, 253.9128, 253.9133, 253.9141, 253.9142, 253.9143, 253.9147, 
    253.915, 253.9144, 253.9151, 253.9124, 253.9138, 253.9116, 253.9123, 
    253.9127, 253.9125, 253.9136, 253.9138, 253.9148, 253.9143, 253.9174, 
    253.916, 253.9198, 253.9187, 253.9116, 253.912, 253.9131, 253.9126, 
    253.9142, 253.9145, 253.9149, 253.9153, 253.9153, 253.9155, 253.9152, 
    253.9155, 253.9141, 253.9147, 253.913, 253.9134, 253.9132, 253.913, 
    253.9137, 253.9144, 253.9144, 253.9146, 253.9152, 253.9142, 253.9175, 
    253.9154, 253.9123, 253.9129, 253.9131, 253.9128, 253.9145, 253.9139, 
    253.9155, 253.9151, 253.9158, 253.9155, 253.9154, 253.9149, 253.9147, 
    253.9139, 253.9133, 253.9129, 253.913, 253.9135, 253.9144, 253.9153, 
    253.9151, 253.9158, 253.914, 253.9148, 253.9145, 253.9152, 253.9136, 
    253.9149, 253.9133, 253.9134, 253.9139, 253.9148, 253.915, 253.9152, 
    253.9151, 253.9144, 253.9143, 253.9139, 253.9137, 253.9134, 253.9131, 
    253.9134, 253.9136, 253.9144, 253.9152, 253.916, 253.9162, 253.9171, 
    253.9163, 253.9175, 253.9164, 253.9183, 253.915, 253.9164, 253.9139, 
    253.9142, 253.9147, 253.9158, 253.9152, 253.9159, 253.9143, 253.9135, 
    253.9133, 253.9129, 253.9133, 253.9133, 253.9137, 253.9135, 253.9145, 
    253.914, 253.9154, 253.9159, 253.9174, 253.9183, 253.9193, 253.9197, 
    253.9198, 253.9199 ;

 TWS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 T_SCALAR =
  0.1456411, 0.1456402, 0.1456404, 0.1456397, 0.1456401, 0.1456396, 
    0.1456409, 0.1456402, 0.1456406, 0.145641, 0.1456385, 0.1456397, 
    0.1456373, 0.145638, 0.1456362, 0.1456374, 0.145636, 0.1456362, 
    0.1456355, 0.1456357, 0.1456349, 0.1456354, 0.1456345, 0.145635, 
    0.1456349, 0.1456355, 0.1456394, 0.1456386, 0.1456395, 0.1456393, 
    0.1456394, 0.1456401, 0.1456404, 0.1456411, 0.145641, 0.1456405, 
    0.1456393, 0.1456397, 0.1456387, 0.1456387, 0.1456377, 0.1456382, 
    0.1456365, 0.145637, 0.1456357, 0.145636, 0.1456357, 0.1456358, 
    0.1456357, 0.1456362, 0.145636, 0.1456364, 0.1456381, 0.1456376, 
    0.1456392, 0.1456402, 0.1456409, 0.1456414, 0.1456413, 0.1456412, 
    0.1456405, 0.1456398, 0.1456393, 0.145639, 0.1456387, 0.1456379, 
    0.1456374, 0.1456364, 0.1456366, 0.1456363, 0.145636, 0.1456356, 
    0.1456357, 0.1456355, 0.1456363, 0.1456358, 0.1456367, 0.1456364, 
    0.1456387, 0.1456396, 0.14564, 0.1456403, 0.1456412, 0.1456406, 
    0.1456409, 0.1456403, 0.1456399, 0.1456401, 0.145639, 0.1456394, 
    0.1456374, 0.1456382, 0.1456361, 0.1456365, 0.145636, 0.1456362, 
    0.1456358, 0.1456362, 0.1456354, 0.1456353, 0.1456354, 0.145635, 
    0.1456362, 0.1456357, 0.1456401, 0.1456401, 0.1456399, 0.1456405, 
    0.1456406, 0.1456411, 0.1456406, 0.1456404, 0.1456399, 0.1456396, 
    0.1456393, 0.1456387, 0.145638, 0.1456372, 0.1456365, 0.1456361, 
    0.1456364, 0.1456362, 0.1456364, 0.1456365, 0.1456353, 0.145636, 
    0.145635, 0.1456351, 0.1456355, 0.1456351, 0.1456401, 0.1456402, 
    0.1456408, 0.1456403, 0.1456412, 0.1456407, 0.1456404, 0.1456394, 
    0.1456392, 0.145639, 0.1456386, 0.1456381, 0.1456373, 0.1456366, 
    0.145636, 0.1456361, 0.1456361, 0.1456359, 0.1456362, 0.1456359, 
    0.1456358, 0.145636, 0.1456351, 0.1456353, 0.1456351, 0.1456352, 
    0.1456402, 0.1456399, 0.14564, 0.1456398, 0.14564, 0.1456391, 0.1456388, 
    0.1456377, 0.1456382, 0.1456374, 0.1456381, 0.145638, 0.1456374, 
    0.145638, 0.1456366, 0.1456376, 0.1456359, 0.1456368, 0.1456359, 
    0.145636, 0.1456358, 0.1456355, 0.1456353, 0.1456348, 0.1456349, 
    0.1456345, 0.1456395, 0.1456391, 0.1456392, 0.1456388, 0.1456385, 
    0.145638, 0.1456371, 0.1456374, 0.1456369, 0.1456368, 0.1456376, 
    0.1456371, 0.1456389, 0.1456386, 0.1456388, 0.1456394, 0.1456374, 
    0.1456384, 0.1456365, 0.1456371, 0.1456356, 0.1456363, 0.1456349, 
    0.1456345, 0.145634, 0.1456336, 0.1456389, 0.1456392, 0.1456387, 
    0.1456382, 0.1456377, 0.145637, 0.145637, 0.1456368, 0.1456365, 
    0.1456363, 0.1456368, 0.1456362, 0.1456385, 0.1456373, 0.1456393, 
    0.1456386, 0.1456382, 0.1456384, 0.1456375, 0.1456373, 0.1456364, 
    0.1456369, 0.1456346, 0.1456355, 0.1456332, 0.1456338, 0.1456393, 
    0.1456389, 0.1456379, 0.1456384, 0.145637, 0.1456366, 0.1456364, 
    0.1456361, 0.145636, 0.1456358, 0.1456361, 0.1456359, 0.145637, 
    0.1456365, 0.145638, 0.1456376, 0.1456378, 0.145638, 0.1456374, 
    0.1456368, 0.1456368, 0.1456366, 0.1456361, 0.145637, 0.1456345, 
    0.1456359, 0.1456386, 0.145638, 0.1456379, 0.1456382, 0.1456367, 
    0.1456372, 0.1456358, 0.1456362, 0.1456356, 0.1456359, 0.1456359, 
    0.1456363, 0.1456365, 0.1456372, 0.1456377, 0.1456381, 0.145638, 
    0.1456376, 0.1456368, 0.145636, 0.1456362, 0.1456357, 0.1456371, 
    0.1456365, 0.1456367, 0.1456361, 0.1456374, 0.1456363, 0.1456378, 
    0.1456376, 0.1456372, 0.1456364, 0.1456362, 0.1456361, 0.1456362, 
    0.1456367, 0.1456368, 0.1456372, 0.1456373, 0.1456376, 0.1456379, 
    0.1456377, 0.1456374, 0.1456367, 0.1456361, 0.1456355, 0.1456354, 
    0.1456348, 0.1456353, 0.1456345, 0.1456351, 0.145634, 0.1456362, 
    0.1456352, 0.1456372, 0.145637, 0.1456365, 0.1456356, 0.1456361, 
    0.1456356, 0.1456368, 0.1456375, 0.1456377, 0.1456381, 0.1456377, 
    0.1456378, 0.1456374, 0.1456375, 0.1456367, 0.1456371, 0.1456359, 
    0.1456356, 0.1456345, 0.145634, 0.1456335, 0.1456333, 0.1456332, 0.1456332,
  0.1512731, 0.1512778, 0.1512769, 0.1512807, 0.1512786, 0.1512811, 
    0.1512741, 0.151278, 0.1512755, 0.1512736, 0.151288, 0.1512809, 
    0.1512957, 0.1512911, 0.1513027, 0.1512949, 0.1513043, 0.1513026, 
    0.1513081, 0.1513065, 0.1513134, 0.1513088, 0.1513171, 0.1513123, 
    0.1513131, 0.1513086, 0.1512824, 0.151287, 0.1512821, 0.1512828, 
    0.1512825, 0.1512786, 0.1512767, 0.1512728, 0.1512735, 0.1512764, 
    0.1512831, 0.1512809, 0.1512866, 0.1512865, 0.1512928, 0.1512899, 
    0.1513007, 0.1512977, 0.1513066, 0.1513043, 0.1513065, 0.1513058, 
    0.1513065, 0.1513031, 0.1513046, 0.1513017, 0.1512904, 0.1512937, 
    0.151284, 0.151278, 0.1512742, 0.1512715, 0.1512719, 0.1512726, 
    0.1512764, 0.15128, 0.1512828, 0.1512846, 0.1512864, 0.1512917, 
    0.1512947, 0.1513013, 0.1513001, 0.1513021, 0.1513041, 0.1513073, 
    0.1513068, 0.1513082, 0.1513021, 0.1513061, 0.1512995, 0.1513013, 
    0.1512866, 0.1512814, 0.151279, 0.1512771, 0.1512722, 0.1512756, 
    0.1512742, 0.1512775, 0.1512795, 0.1512785, 0.1512847, 0.1512823, 
    0.1512949, 0.1512894, 0.1513039, 0.1513004, 0.1513047, 0.1513025, 
    0.1513062, 0.1513029, 0.1513088, 0.15131, 0.1513091, 0.1513126, 
    0.1513027, 0.1513064, 0.1512784, 0.1512786, 0.1512794, 0.151276, 
    0.1512758, 0.1512728, 0.1512755, 0.1512766, 0.1512796, 0.1512813, 
    0.151283, 0.1512866, 0.1512907, 0.1512964, 0.1513006, 0.1513034, 
    0.1513017, 0.1513032, 0.1513015, 0.1513007, 0.1513095, 0.1513046, 
    0.1513121, 0.1513117, 0.1513082, 0.1513117, 0.1512787, 0.1512778, 
    0.1512745, 0.1512771, 0.1512724, 0.151275, 0.1512765, 0.1512822, 
    0.1512836, 0.1512847, 0.1512871, 0.1512901, 0.1512953, 0.1512999, 
    0.1513042, 0.1513039, 0.151304, 0.1513049, 0.1513026, 0.1513053, 
    0.1513058, 0.1513046, 0.1513116, 0.1513096, 0.1513117, 0.1513103, 
    0.1512781, 0.1512797, 0.1512788, 0.1512804, 0.1512793, 0.1512842, 
    0.1512858, 0.1512929, 0.15129, 0.1512946, 0.1512905, 0.1512912, 
    0.1512946, 0.1512907, 0.1512996, 0.1512935, 0.151305, 0.1512987, 
    0.1513054, 0.1513042, 0.1513062, 0.1513079, 0.1513101, 0.1513142, 
    0.1513133, 0.1513168, 0.151282, 0.151284, 0.1512839, 0.1512861, 
    0.1512876, 0.1512911, 0.1512967, 0.1512946, 0.1512984, 0.1512992, 
    0.1512934, 0.1512969, 0.1512854, 0.1512872, 0.1512862, 0.1512822, 
    0.151295, 0.1512884, 0.1513007, 0.1512971, 0.1513077, 0.1513023, 
    0.1513128, 0.1513171, 0.1513215, 0.1513264, 0.1512852, 0.1512838, 
    0.1512863, 0.1512897, 0.151293, 0.1512973, 0.1512978, 0.1512986, 
    0.1513007, 0.1513024, 0.1512988, 0.1513029, 0.1512875, 0.1512956, 
    0.1512832, 0.1512869, 0.1512895, 0.1512884, 0.1512944, 0.1512958, 
    0.1513014, 0.1512985, 0.151316, 0.1513082, 0.1513303, 0.151324, 
    0.1512833, 0.1512852, 0.1512917, 0.1512886, 0.1512976, 0.1512998, 
    0.1513016, 0.1513039, 0.1513042, 0.1513055, 0.1513033, 0.1513055, 
    0.1512973, 0.1513009, 0.151291, 0.1512934, 0.1512923, 0.1512911, 
    0.1512949, 0.1512988, 0.151299, 0.1513002, 0.1513036, 0.1512976, 
    0.1513169, 0.1513048, 0.1512873, 0.1512908, 0.1512914, 0.15129, 
    0.1512996, 0.1512961, 0.1513055, 0.151303, 0.1513072, 0.1513051, 
    0.1513048, 0.1513021, 0.1513004, 0.1512962, 0.1512929, 0.1512902, 
    0.1512908, 0.1512937, 0.1512991, 0.1513042, 0.151303, 0.1513069, 
    0.1512969, 0.151301, 0.1512994, 0.1513036, 0.1512945, 0.151302, 
    0.1512926, 0.1512934, 0.151296, 0.1513012, 0.1513025, 0.1513038, 
    0.151303, 0.1512992, 0.1512986, 0.151296, 0.1512952, 0.1512932, 
    0.1512916, 0.1512931, 0.1512946, 0.1512993, 0.1513034, 0.1513079, 
    0.1513091, 0.1513142, 0.1513099, 0.1513169, 0.1513108, 0.1513215, 
    0.1513026, 0.1513108, 0.1512962, 0.1512978, 0.1513005, 0.1513071, 
    0.1513036, 0.1513077, 0.1512986, 0.1512938, 0.1512927, 0.1512904, 
    0.1512927, 0.1512925, 0.1512948, 0.1512941, 0.1512994, 0.1512965, 
    0.1513047, 0.1513077, 0.1513164, 0.1513217, 0.1513272, 0.1513296, 
    0.1513304, 0.1513307,
  0.1611241, 0.1611301, 0.1611289, 0.1611337, 0.1611311, 0.1611342, 
    0.1611253, 0.1611303, 0.1611271, 0.1611246, 0.161143, 0.1611339, 
    0.1611529, 0.161147, 0.1611619, 0.1611519, 0.161164, 0.1611618, 
    0.1611688, 0.1611668, 0.1611757, 0.1611697, 0.1611805, 0.1611743, 
    0.1611752, 0.1611695, 0.1611359, 0.1611418, 0.1611355, 0.1611363, 
    0.161136, 0.1611311, 0.1611286, 0.1611236, 0.1611246, 0.1611282, 
    0.1611367, 0.1611339, 0.1611412, 0.1611411, 0.1611492, 0.1611455, 
    0.1611593, 0.1611554, 0.1611669, 0.161164, 0.1611667, 0.1611659, 
    0.1611667, 0.1611625, 0.1611643, 0.1611606, 0.1611462, 0.1611504, 
    0.1611379, 0.1611303, 0.1611255, 0.1611221, 0.1611225, 0.1611235, 
    0.1611283, 0.1611329, 0.1611364, 0.1611387, 0.161141, 0.1611478, 
    0.1611516, 0.1611601, 0.1611586, 0.1611611, 0.1611637, 0.1611678, 
    0.1611671, 0.161169, 0.1611611, 0.1611663, 0.1611578, 0.1611601, 
    0.1611413, 0.1611347, 0.1611316, 0.1611291, 0.1611229, 0.1611272, 
    0.1611255, 0.1611296, 0.1611321, 0.1611309, 0.1611388, 0.1611357, 
    0.1611519, 0.1611449, 0.1611634, 0.1611589, 0.1611645, 0.1611616, 
    0.1611664, 0.1611621, 0.1611697, 0.1611713, 0.1611702, 0.1611746, 
    0.1611619, 0.1611667, 0.1611308, 0.161131, 0.161132, 0.1611277, 
    0.1611275, 0.1611236, 0.1611271, 0.1611285, 0.1611323, 0.1611345, 
    0.1611366, 0.1611413, 0.1611465, 0.1611538, 0.1611592, 0.1611628, 
    0.1611606, 0.1611626, 0.1611604, 0.1611594, 0.1611707, 0.1611643, 
    0.1611739, 0.1611734, 0.161169, 0.1611735, 0.1611312, 0.16113, 0.1611258, 
    0.1611291, 0.1611232, 0.1611265, 0.1611283, 0.1611357, 0.1611374, 
    0.1611389, 0.1611419, 0.1611457, 0.1611524, 0.1611583, 0.1611638, 
    0.1611634, 0.1611636, 0.1611648, 0.1611618, 0.1611653, 0.1611658, 
    0.1611643, 0.1611733, 0.1611708, 0.1611734, 0.1611717, 0.1611304, 
    0.1611324, 0.1611313, 0.1611333, 0.1611319, 0.1611383, 0.1611402, 
    0.1611492, 0.1611456, 0.1611515, 0.1611462, 0.1611471, 0.1611516, 
    0.1611465, 0.1611579, 0.1611501, 0.1611648, 0.1611568, 0.1611653, 
    0.1611638, 0.1611663, 0.1611686, 0.1611715, 0.1611767, 0.1611755, 
    0.16118, 0.1611354, 0.161138, 0.1611378, 0.1611406, 0.1611426, 0.161147, 
    0.1611541, 0.1611515, 0.1611564, 0.1611574, 0.1611499, 0.1611544, 
    0.1611398, 0.1611421, 0.1611407, 0.1611356, 0.161152, 0.1611435, 
    0.1611593, 0.1611547, 0.1611682, 0.1611614, 0.1611748, 0.1611805, 
    0.1611861, 0.1611924, 0.1611395, 0.1611377, 0.1611409, 0.1611452, 
    0.1611494, 0.1611549, 0.1611555, 0.1611566, 0.1611593, 0.1611615, 
    0.1611568, 0.1611621, 0.1611425, 0.1611528, 0.161137, 0.1611416, 
    0.161145, 0.1611436, 0.1611512, 0.161153, 0.1611602, 0.1611565, 0.161179, 
    0.161169, 0.1611974, 0.1611893, 0.1611371, 0.1611395, 0.1611478, 
    0.1611438, 0.1611553, 0.1611582, 0.1611605, 0.1611634, 0.1611638, 
    0.1611655, 0.1611627, 0.1611654, 0.161155, 0.1611596, 0.1611469, 0.16115, 
    0.1611486, 0.161147, 0.1611518, 0.1611569, 0.1611571, 0.1611587, 
    0.161163, 0.1611554, 0.1611801, 0.1611646, 0.1611421, 0.1611466, 
    0.1611474, 0.1611456, 0.1611579, 0.1611534, 0.1611655, 0.1611622, 
    0.1611676, 0.1611649, 0.1611645, 0.1611611, 0.161159, 0.1611536, 
    0.1611492, 0.1611459, 0.1611467, 0.1611504, 0.1611572, 0.1611638, 
    0.1611623, 0.1611672, 0.1611545, 0.1611598, 0.1611577, 0.1611631, 
    0.1611514, 0.1611611, 0.1611489, 0.16115, 0.1611533, 0.16116, 0.1611617, 
    0.1611633, 0.1611623, 0.1611574, 0.1611566, 0.1611533, 0.1611523, 
    0.1611497, 0.1611476, 0.1611495, 0.1611515, 0.1611574, 0.1611627, 
    0.1611686, 0.1611701, 0.1611767, 0.1611712, 0.1611802, 0.1611723, 
    0.1611861, 0.1611618, 0.1611723, 0.1611535, 0.1611555, 0.1611591, 
    0.1611676, 0.1611631, 0.1611684, 0.1611566, 0.1611505, 0.161149, 
    0.1611461, 0.1611491, 0.1611488, 0.1611517, 0.1611508, 0.1611577, 
    0.161154, 0.1611645, 0.1611684, 0.1611795, 0.1611863, 0.1611934, 
    0.1611966, 0.1611975, 0.1611979,
  0.175334, 0.1753385, 0.1753377, 0.1753413, 0.1753393, 0.1753417, 0.175335, 
    0.1753387, 0.1753363, 0.1753345, 0.1753483, 0.1753415, 0.1753558, 
    0.1753513, 0.1753628, 0.1753551, 0.1753644, 0.1753627, 0.1753681, 
    0.1753666, 0.1753735, 0.1753689, 0.1753772, 0.1753724, 0.1753731, 
    0.1753687, 0.1753429, 0.1753474, 0.1753426, 0.1753433, 0.175343, 
    0.1753393, 0.1753374, 0.1753338, 0.1753344, 0.1753372, 0.1753436, 
    0.1753414, 0.175347, 0.1753468, 0.175353, 0.1753502, 0.1753608, 
    0.1753578, 0.1753667, 0.1753644, 0.1753665, 0.1753659, 0.1753665, 
    0.1753632, 0.1753646, 0.1753618, 0.1753507, 0.1753539, 0.1753444, 
    0.1753387, 0.1753351, 0.1753326, 0.1753329, 0.1753336, 0.1753372, 
    0.1753407, 0.1753433, 0.1753451, 0.1753468, 0.175352, 0.1753549, 
    0.1753614, 0.1753603, 0.1753622, 0.1753642, 0.1753674, 0.1753669, 
    0.1753683, 0.1753622, 0.1753662, 0.1753596, 0.1753614, 0.175347, 
    0.175342, 0.1753397, 0.1753378, 0.1753332, 0.1753364, 0.1753351, 
    0.1753382, 0.1753401, 0.1753392, 0.1753451, 0.1753428, 0.1753551, 
    0.1753497, 0.1753639, 0.1753605, 0.1753648, 0.1753626, 0.1753663, 
    0.175363, 0.1753688, 0.1753701, 0.1753692, 0.1753726, 0.1753628, 
    0.1753665, 0.1753391, 0.1753393, 0.17534, 0.1753368, 0.1753366, 
    0.1753337, 0.1753363, 0.1753374, 0.1753403, 0.1753419, 0.1753435, 
    0.175347, 0.1753509, 0.1753566, 0.1753607, 0.1753635, 0.1753618, 
    0.1753633, 0.1753616, 0.1753609, 0.1753696, 0.1753646, 0.1753721, 
    0.1753717, 0.1753683, 0.1753718, 0.1753394, 0.1753385, 0.1753354, 
    0.1753378, 0.1753334, 0.1753359, 0.1753372, 0.1753428, 0.1753441, 
    0.1753452, 0.1753475, 0.1753504, 0.1753555, 0.1753601, 0.1753643, 
    0.175364, 0.1753641, 0.175365, 0.1753627, 0.1753654, 0.1753658, 
    0.1753647, 0.1753717, 0.1753697, 0.1753717, 0.1753704, 0.1753388, 
    0.1753403, 0.1753395, 0.175341, 0.1753399, 0.1753447, 0.1753462, 
    0.1753531, 0.1753503, 0.1753548, 0.1753508, 0.1753515, 0.1753549, 
    0.175351, 0.1753597, 0.1753537, 0.1753651, 0.1753588, 0.1753654, 
    0.1753643, 0.1753662, 0.175368, 0.1753702, 0.1753743, 0.1753734, 
    0.1753769, 0.1753426, 0.1753445, 0.1753444, 0.1753465, 0.175348, 
    0.1753514, 0.1753568, 0.1753548, 0.1753586, 0.1753593, 0.1753536, 
    0.1753571, 0.1753459, 0.1753476, 0.1753466, 0.1753427, 0.1753552, 
    0.1753487, 0.1753608, 0.1753572, 0.1753677, 0.1753624, 0.1753728, 
    0.1753773, 0.1753817, 0.1753867, 0.1753456, 0.1753443, 0.1753467, 
    0.17535, 0.1753532, 0.1753574, 0.1753579, 0.1753587, 0.1753608, 
    0.1753625, 0.1753589, 0.175363, 0.1753479, 0.1753558, 0.1753438, 
    0.1753473, 0.1753498, 0.1753488, 0.1753546, 0.1753559, 0.1753615, 
    0.1753586, 0.1753761, 0.1753683, 0.1753906, 0.1753842, 0.1753438, 
    0.1753456, 0.175352, 0.175349, 0.1753577, 0.1753599, 0.1753617, 0.175364, 
    0.1753643, 0.1753656, 0.1753634, 0.1753656, 0.1753574, 0.1753611, 
    0.1753513, 0.1753536, 0.1753526, 0.1753514, 0.175355, 0.1753589, 
    0.1753591, 0.1753603, 0.1753637, 0.1753578, 0.175377, 0.1753649, 
    0.1753476, 0.1753511, 0.1753516, 0.1753503, 0.1753597, 0.1753563, 
    0.1753656, 0.1753631, 0.1753672, 0.1753651, 0.1753648, 0.1753622, 
    0.1753605, 0.1753564, 0.1753531, 0.1753505, 0.1753511, 0.1753539, 
    0.1753592, 0.1753643, 0.1753631, 0.1753669, 0.1753571, 0.1753611, 
    0.1753595, 0.1753637, 0.1753547, 0.1753621, 0.1753528, 0.1753536, 
    0.1753562, 0.1753614, 0.1753626, 0.1753639, 0.1753631, 0.1753593, 
    0.1753587, 0.1753561, 0.1753554, 0.1753535, 0.1753518, 0.1753533, 
    0.1753548, 0.1753594, 0.1753635, 0.175368, 0.1753691, 0.1753743, 0.17537, 
    0.1753771, 0.1753709, 0.1753817, 0.1753627, 0.1753709, 0.1753563, 
    0.1753579, 0.1753606, 0.1753672, 0.1753637, 0.1753678, 0.1753587, 
    0.175354, 0.1753529, 0.1753507, 0.1753529, 0.1753528, 0.1753549, 
    0.1753542, 0.1753595, 0.1753567, 0.1753648, 0.1753678, 0.1753765, 
    0.1753818, 0.1753875, 0.17539, 0.1753907, 0.175391,
  0.1899463, 0.1899477, 0.1899474, 0.1899485, 0.1899479, 0.1899486, 
    0.1899466, 0.1899477, 0.189947, 0.1899464, 0.1899507, 0.1899486, 
    0.1899532, 0.1899517, 0.1899556, 0.189953, 0.1899561, 0.1899555, 
    0.1899574, 0.1899568, 0.1899593, 0.1899576, 0.1899606, 0.1899589, 
    0.1899591, 0.1899576, 0.189949, 0.1899505, 0.1899489, 0.1899491, 
    0.1899491, 0.1899479, 0.1899473, 0.1899462, 0.1899464, 0.1899472, 
    0.1899492, 0.1899486, 0.1899503, 0.1899503, 0.1899523, 0.1899514, 
    0.1899549, 0.1899539, 0.1899569, 0.1899561, 0.1899568, 0.1899566, 
    0.1899568, 0.1899557, 0.1899562, 0.1899552, 0.1899515, 0.1899526, 
    0.1899495, 0.1899477, 0.1899466, 0.1899458, 0.189946, 0.1899462, 
    0.1899472, 0.1899483, 0.1899492, 0.1899497, 0.1899503, 0.1899519, 
    0.1899529, 0.1899551, 0.1899547, 0.1899554, 0.189956, 0.1899571, 
    0.1899569, 0.1899574, 0.1899554, 0.1899567, 0.1899545, 0.1899551, 
    0.1899503, 0.1899488, 0.189948, 0.1899475, 0.189946, 0.189947, 0.1899466, 
    0.1899476, 0.1899482, 0.1899479, 0.1899497, 0.189949, 0.189953, 
    0.1899512, 0.1899559, 0.1899548, 0.1899562, 0.1899555, 0.1899568, 
    0.1899556, 0.1899576, 0.1899581, 0.1899578, 0.189959, 0.1899555, 
    0.1899568, 0.1899479, 0.1899479, 0.1899481, 0.1899471, 0.1899471, 
    0.1899462, 0.189947, 0.1899473, 0.1899482, 0.1899487, 0.1899492, 
    0.1899503, 0.1899516, 0.1899535, 0.1899548, 0.1899558, 0.1899552, 
    0.1899557, 0.1899552, 0.1899549, 0.1899579, 0.1899562, 0.1899588, 
    0.1899586, 0.1899574, 0.1899587, 0.1899479, 0.1899477, 0.1899467, 
    0.1899475, 0.1899461, 0.1899468, 0.1899473, 0.189949, 0.1899494, 
    0.1899498, 0.1899505, 0.1899514, 0.1899531, 0.1899546, 0.1899561, 
    0.189956, 0.189956, 0.1899563, 0.1899555, 0.1899564, 0.1899566, 
    0.1899562, 0.1899586, 0.1899579, 0.1899586, 0.1899582, 0.1899478, 
    0.1899482, 0.189948, 0.1899484, 0.1899481, 0.1899496, 0.1899501, 
    0.1899523, 0.1899514, 0.1899529, 0.1899515, 0.1899518, 0.1899529, 
    0.1899516, 0.1899545, 0.1899525, 0.1899563, 0.1899542, 0.1899565, 
    0.1899561, 0.1899567, 0.1899573, 0.1899581, 0.1899596, 0.1899592, 
    0.1899605, 0.1899489, 0.1899495, 0.1899495, 0.1899502, 0.1899506, 
    0.1899517, 0.1899535, 0.1899529, 0.1899541, 0.1899544, 0.1899525, 
    0.1899536, 0.18995, 0.1899505, 0.1899502, 0.189949, 0.189953, 0.1899509, 
    0.1899549, 0.1899537, 0.1899572, 0.1899554, 0.189959, 0.1899606, 
    0.1899622, 0.189964, 0.1899499, 0.1899495, 0.1899502, 0.1899513, 
    0.1899523, 0.1899537, 0.1899539, 0.1899542, 0.1899549, 0.1899555, 
    0.1899542, 0.1899556, 0.1899506, 0.1899532, 0.1899493, 0.1899504, 
    0.1899512, 0.1899509, 0.1899528, 0.1899532, 0.1899551, 0.1899541, 
    0.1899602, 0.1899574, 0.1899655, 0.1899631, 0.1899493, 0.1899499, 
    0.1899519, 0.189951, 0.1899538, 0.1899546, 0.1899552, 0.1899559, 
    0.1899561, 0.1899565, 0.1899558, 0.1899565, 0.1899537, 0.189955, 
    0.1899517, 0.1899525, 0.1899521, 0.1899517, 0.189953, 0.1899542, 
    0.1899543, 0.1899547, 0.1899558, 0.1899539, 0.1899605, 0.1899563, 
    0.1899505, 0.1899516, 0.1899518, 0.1899514, 0.1899545, 0.1899533, 
    0.1899565, 0.1899556, 0.1899571, 0.1899564, 0.1899562, 0.1899554, 
    0.1899548, 0.1899534, 0.1899523, 0.1899515, 0.1899517, 0.1899526, 
    0.1899543, 0.1899561, 0.1899557, 0.189957, 0.1899536, 0.189955, 
    0.1899544, 0.1899559, 0.1899528, 0.1899553, 0.1899522, 0.1899525, 
    0.1899533, 0.1899551, 0.1899555, 0.1899559, 0.1899557, 0.1899544, 
    0.1899542, 0.1899533, 0.1899531, 0.1899524, 0.1899519, 0.1899524, 
    0.1899529, 0.1899544, 0.1899558, 0.1899573, 0.1899577, 0.1899596, 
    0.189958, 0.1899605, 0.1899583, 0.1899622, 0.1899555, 0.1899583, 
    0.1899534, 0.1899539, 0.1899548, 0.1899571, 0.1899559, 0.1899573, 
    0.1899542, 0.1899526, 0.1899522, 0.1899515, 0.1899523, 0.1899522, 
    0.1899529, 0.1899527, 0.1899544, 0.1899535, 0.1899562, 0.1899573, 
    0.1899603, 0.1899623, 0.1899643, 0.1899652, 0.1899655, 0.1899657,
  0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973189, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973188, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.197319, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973189, 0.1973189, 0.197319, 0.197319, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973188, 0.1973189, 0.1973188, 0.1973188, 
    0.1973188, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973189, 
    0.1973188, 0.1973188, 0.1973189, 0.1973188, 0.1973189, 0.1973188, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973188, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 
    0.1973188, 0.1973189, 0.1973188, 0.1973188, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973188, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973188, 
    0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.197319, 
    0.1973189, 0.197319, 0.1973189, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973188, 
    0.1973189, 0.197319, 0.1973191, 0.1973192, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.197319, 0.1973189, 0.1973192, 0.1973191, 
    0.1973189, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973188, 
    0.197319, 0.1973189, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973189, 0.1973189, 0.1973189, 0.1973189, 
    0.1973189, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973189, 0.1973189, 
    0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 
    0.1973189, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 0.1973189, 
    0.1973189, 0.197319, 0.1973189, 0.197319, 0.1973189, 0.1973191, 
    0.1973188, 0.1973189, 0.1973188, 0.1973188, 0.1973188, 0.1973189, 
    0.1973189, 0.1973189, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 0.1973188, 
    0.1973189, 0.1973189, 0.197319, 0.1973191, 0.1973192, 0.1973192, 
    0.1973192, 0.1973193,
  0.1984799, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984799, 0.1984798, 0.1984799, 0.1984799, 0.1984798, 0.1984798, 
    0.1984797, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984799, 0.1984799, 0.1984799, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984799, 0.1984799, 0.1984799, 0.1984799, 
    0.1984799, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984799, 0.1984799, 
    0.1984799, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984799, 
    0.1984799, 0.1984799, 0.1984799, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 
    0.1984799, 0.1984798, 0.1984799, 0.1984799, 0.1984799, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984798, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984798, 0.1984797, 0.1984797, 
    0.1984798, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984797, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984796, 0.1984796, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984797, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984796, 0.1984796, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 0.1984798, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984797, 
    0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984796, 
    0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984798, 0.1984798, 0.1984798, 
    0.1984798, 0.1984798, 0.1984798, 0.1984798, 0.1984797, 0.1984797, 
    0.1984797, 0.1984797, 0.1984797, 0.1984796, 0.1984796, 0.1984796, 
    0.1984796, 0.1984796,
  0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 U10 =
  5.611711, 5.611763, 5.611753, 5.611795, 5.611772, 5.611799, 5.611722, 
    5.611765, 5.611738, 5.611716, 5.611874, 5.611797, 5.611958, 5.611908, 
    5.612037, 5.61195, 5.612055, 5.612035, 5.612096, 5.612079, 5.612154, 
    5.612104, 5.612195, 5.612143, 5.612151, 5.612103, 5.611814, 5.611864, 
    5.61181, 5.611817, 5.611814, 5.611773, 5.61175, 5.611707, 5.611715, 
    5.611747, 5.611821, 5.611797, 5.61186, 5.611858, 5.611928, 5.611896, 
    5.612014, 5.61198, 5.61208, 5.612055, 5.612079, 5.612072, 5.612079, 
    5.612041, 5.612058, 5.612025, 5.611902, 5.611937, 5.611831, 5.611764, 
    5.611723, 5.611693, 5.611698, 5.611705, 5.611747, 5.611788, 5.611818, 
    5.611838, 5.611858, 5.611915, 5.611948, 5.61202, 5.612008, 5.61203, 
    5.612052, 5.612088, 5.612082, 5.612098, 5.61203, 5.612075, 5.612, 
    5.612021, 5.611859, 5.611804, 5.611776, 5.611755, 5.611701, 5.611738, 
    5.611723, 5.611759, 5.611782, 5.611771, 5.611839, 5.611812, 5.611949, 
    5.611891, 5.61205, 5.61201, 5.612059, 5.612035, 5.612076, 5.612039, 
    5.612104, 5.612117, 5.612108, 5.612145, 5.612037, 5.612078, 5.61177, 
    5.611772, 5.611781, 5.611742, 5.611741, 5.611707, 5.611737, 5.61175, 
    5.611783, 5.611802, 5.61182, 5.61186, 5.611904, 5.611967, 5.612013, 
    5.612045, 5.612026, 5.612042, 5.612023, 5.612015, 5.612112, 5.612057, 
    5.61214, 5.612136, 5.612098, 5.612136, 5.611773, 5.611763, 5.611726, 
    5.611755, 5.611703, 5.611732, 5.611748, 5.611812, 5.611827, 5.611839, 
    5.611866, 5.611898, 5.611955, 5.612005, 5.612054, 5.61205, 5.612051, 
    5.612062, 5.612036, 5.612066, 5.612071, 5.612058, 5.612135, 5.612113, 
    5.612135, 5.612122, 5.611766, 5.611784, 5.611774, 5.611792, 5.611779, 
    5.611834, 5.61185, 5.611928, 5.611897, 5.611947, 5.611902, 5.61191, 
    5.611947, 5.611905, 5.612001, 5.611934, 5.612062, 5.61199, 5.612067, 
    5.612053, 5.612075, 5.612094, 5.612119, 5.612164, 5.612154, 5.612191, 
    5.61181, 5.611832, 5.611831, 5.611854, 5.611871, 5.611909, 5.611969, 
    5.611947, 5.611989, 5.611997, 5.611934, 5.611971, 5.611847, 5.611866, 
    5.611856, 5.611811, 5.611951, 5.611879, 5.612013, 5.611974, 5.612092, 
    5.612032, 5.612148, 5.612195, 5.612242, 5.612293, 5.611845, 5.61183, 
    5.611857, 5.611894, 5.611929, 5.611976, 5.611981, 5.611989, 5.612013, 
    5.612034, 5.611991, 5.612039, 5.611869, 5.611958, 5.611823, 5.611863, 
    5.611892, 5.61188, 5.611944, 5.611959, 5.612021, 5.611989, 5.612182, 
    5.612097, 5.612335, 5.612268, 5.611824, 5.611845, 5.611916, 5.611882, 
    5.611979, 5.612003, 5.612025, 5.61205, 5.612053, 5.612068, 5.612044, 
    5.612068, 5.611976, 5.612017, 5.611908, 5.611934, 5.611922, 5.611909, 
    5.61195, 5.611992, 5.611994, 5.612008, 5.612045, 5.61198, 5.612191, 
    5.612059, 5.611867, 5.611905, 5.611912, 5.611897, 5.612, 5.611963, 
    5.612068, 5.61204, 5.612086, 5.612063, 5.61206, 5.61203, 5.612011, 
    5.611965, 5.611928, 5.611899, 5.611906, 5.611938, 5.611995, 5.612053, 
    5.61204, 5.612083, 5.611972, 5.612018, 5.611999, 5.612047, 5.611946, 
    5.612028, 5.611925, 5.611934, 5.611962, 5.61202, 5.612035, 5.612049, 
    5.612041, 5.611996, 5.61199, 5.611962, 5.611953, 5.611932, 5.611914, 
    5.61193, 5.611947, 5.611997, 5.612044, 5.612094, 5.612107, 5.612163, 
    5.612116, 5.612191, 5.612125, 5.612241, 5.612035, 5.612125, 5.611964, 
    5.611981, 5.612011, 5.612085, 5.612047, 5.612092, 5.61199, 5.611938, 
    5.611926, 5.611901, 5.611927, 5.611925, 5.611949, 5.611941, 5.611999, 
    5.611968, 5.61206, 5.612092, 5.612186, 5.612243, 5.612302, 5.612328, 
    5.612336, 5.612339 ;

 URBAN_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 URBAN_HEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 VOCFLXT =
  5.912984e-15, 5.911853e-15, 5.912067e-15, 5.911168e-15, 5.911659e-15, 
    5.911075e-15, 5.912745e-15, 5.911816e-15, 5.912404e-15, 5.912869e-15, 
    5.909452e-15, 5.911124e-15, 5.90763e-15, 5.908707e-15, 5.905975e-15, 
    5.907809e-15, 5.905602e-15, 5.906006e-15, 5.904739e-15, 5.9051e-15, 
    5.903526e-15, 5.904571e-15, 5.902678e-15, 5.903764e-15, 5.903602e-15, 
    5.90461e-15, 5.910767e-15, 5.909667e-15, 5.910838e-15, 5.910679e-15, 
    5.910746e-15, 5.911656e-15, 5.912129e-15, 5.913056e-15, 5.912884e-15, 
    5.912195e-15, 5.910608e-15, 5.911132e-15, 5.90977e-15, 5.909801e-15, 
    5.908301e-15, 5.908977e-15, 5.906447e-15, 5.907161e-15, 5.905085e-15, 
    5.905609e-15, 5.905113e-15, 5.90526e-15, 5.905111e-15, 5.905879e-15, 
    5.905551e-15, 5.90622e-15, 5.908855e-15, 5.908087e-15, 5.910392e-15, 
    5.911814e-15, 5.912708e-15, 5.913359e-15, 5.913267e-15, 5.913096e-15, 
    5.912191e-15, 5.911324e-15, 5.910669e-15, 5.910235e-15, 5.909805e-15, 
    5.908559e-15, 5.907854e-15, 5.906313e-15, 5.906572e-15, 5.906119e-15, 
    5.90566e-15, 5.904915e-15, 5.905035e-15, 5.904711e-15, 5.906118e-15, 
    5.905189e-15, 5.906726e-15, 5.906307e-15, 5.90976e-15, 5.910987e-15, 
    5.911572e-15, 5.912029e-15, 5.913198e-15, 5.912395e-15, 5.912713e-15, 
    5.911941e-15, 5.91146e-15, 5.911695e-15, 5.910223e-15, 5.910797e-15, 
    5.907813e-15, 5.909096e-15, 5.905714e-15, 5.906518e-15, 5.905518e-15, 
    5.906024e-15, 5.905163e-15, 5.905938e-15, 5.904585e-15, 5.904299e-15, 
    5.904496e-15, 5.903716e-15, 5.905983e-15, 5.90512e-15, 5.911705e-15, 
    5.911667e-15, 5.911483e-15, 5.912295e-15, 5.912341e-15, 5.913065e-15, 
    5.912414e-15, 5.912143e-15, 5.911427e-15, 5.911017e-15, 5.910623e-15, 
    5.909757e-15, 5.908802e-15, 5.907449e-15, 5.906467e-15, 5.905813e-15, 
    5.906209e-15, 5.90586e-15, 5.906253e-15, 5.906434e-15, 5.904411e-15, 
    5.905552e-15, 5.903828e-15, 5.90392e-15, 5.904706e-15, 5.90391e-15, 
    5.911639e-15, 5.911859e-15, 5.912646e-15, 5.91203e-15, 5.913143e-15, 
    5.912529e-15, 5.912181e-15, 5.910801e-15, 5.910481e-15, 5.910208e-15, 
    5.90965e-15, 5.908943e-15, 5.90771e-15, 5.906627e-15, 5.905631e-15, 
    5.905702e-15, 5.905678e-15, 5.905462e-15, 5.906005e-15, 5.905373e-15, 
    5.905274e-15, 5.905544e-15, 5.903934e-15, 5.904392e-15, 5.903923e-15, 
    5.904219e-15, 5.911786e-15, 5.911412e-15, 5.911615e-15, 5.911238e-15, 
    5.911509e-15, 5.910324e-15, 5.909969e-15, 5.908291e-15, 5.908961e-15, 
    5.907874e-15, 5.908845e-15, 5.908677e-15, 5.907869e-15, 5.908787e-15, 
    5.9067e-15, 5.908142e-15, 5.905454e-15, 5.906919e-15, 5.905364e-15, 
    5.905635e-15, 5.90518e-15, 5.90478e-15, 5.904264e-15, 5.903335e-15, 
    5.903547e-15, 5.902759e-15, 5.91085e-15, 5.910374e-15, 5.910402e-15, 
    5.909894e-15, 5.909522e-15, 5.908698e-15, 5.907395e-15, 5.90788e-15, 
    5.906975e-15, 5.906798e-15, 5.908166e-15, 5.907339e-15, 5.910044e-15, 
    5.909621e-15, 5.909863e-15, 5.91082e-15, 5.907787e-15, 5.90935e-15, 
    5.906453e-15, 5.907295e-15, 5.904839e-15, 5.906072e-15, 5.903667e-15, 
    5.902677e-15, 5.901684e-15, 5.900599e-15, 5.910099e-15, 5.910424e-15, 
    5.90983e-15, 5.909033e-15, 5.908256e-15, 5.907247e-15, 5.907136e-15, 
    5.906951e-15, 5.906455e-15, 5.906045e-15, 5.906906e-15, 5.905941e-15, 
    5.909549e-15, 5.907646e-15, 5.910559e-15, 5.909699e-15, 5.909074e-15, 
    5.909335e-15, 5.907932e-15, 5.907608e-15, 5.906292e-15, 5.906964e-15, 
    5.902933e-15, 5.904714e-15, 5.89973e-15, 5.901127e-15, 5.910541e-15, 
    5.910094e-15, 5.908558e-15, 5.909286e-15, 5.907172e-15, 5.906658e-15, 
    5.906229e-15, 5.905704e-15, 5.905637e-15, 5.905325e-15, 5.905839e-15, 
    5.90534e-15, 5.907245e-15, 5.90639e-15, 5.908717e-15, 5.908158e-15, 
    5.908411e-15, 5.908698e-15, 5.907814e-15, 5.906896e-15, 5.906854e-15, 
    5.906563e-15, 5.905784e-15, 5.907163e-15, 5.902743e-15, 5.905505e-15, 
    5.909607e-15, 5.908777e-15, 5.908632e-15, 5.908958e-15, 5.906711e-15, 
    5.907527e-15, 5.905329e-15, 5.905918e-15, 5.904949e-15, 5.905432e-15, 
    5.905504e-15, 5.90612e-15, 5.90651e-15, 5.907494e-15, 5.908288e-15, 
    5.908908e-15, 5.908762e-15, 5.908081e-15, 5.906834e-15, 5.905642e-15, 
    5.905905e-15, 5.905022e-15, 5.907326e-15, 5.906369e-15, 5.906747e-15, 
    5.905761e-15, 5.907898e-15, 5.906143e-15, 5.908355e-15, 5.908156e-15, 
    5.907543e-15, 5.906319e-15, 5.906016e-15, 5.905733e-15, 5.905904e-15, 
    5.906799e-15, 5.906936e-15, 5.907553e-15, 5.907734e-15, 5.908198e-15, 
    5.908593e-15, 5.908237e-15, 5.907869e-15, 5.90679e-15, 5.905829e-15, 
    5.904778e-15, 5.904512e-15, 5.90334e-15, 5.904323e-15, 5.902732e-15, 
    5.904129e-15, 5.90169e-15, 5.906009e-15, 5.904127e-15, 5.907508e-15, 
    5.907137e-15, 5.90649e-15, 5.904965e-15, 5.905765e-15, 5.904819e-15, 
    5.906939e-15, 5.908068e-15, 5.908334e-15, 5.908874e-15, 5.908322e-15, 
    5.908366e-15, 5.907838e-15, 5.908007e-15, 5.906753e-15, 5.907425e-15, 
    5.905512e-15, 5.904821e-15, 5.902849e-15, 5.901658e-15, 5.900413e-15, 
    5.899875e-15, 5.89971e-15, 5.899642e-15 ;

 VOLR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WA =
  4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000 ;

 WASTEHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WF =
  7.141488, 7.168028, 7.162865, 7.184313, 7.172412, 7.186463, 7.146866, 
    7.169081, 7.154895, 7.143879, 7.226072, 7.185272, 7.268681, 7.242513, 
    7.308392, 7.264599, 7.317247, 7.307134, 7.337627, 7.328882, 7.367975, 
    7.341666, 7.388316, 7.36169, 7.365847, 7.340798, 7.193476, 7.22098, 
    7.191847, 7.195764, 7.194007, 7.172655, 7.161908, 7.139468, 7.143539, 
    7.160026, 7.197526, 7.184784, 7.216947, 7.216219, 7.252151, 7.235933, 
    7.296537, 7.279277, 7.329247, 7.316654, 7.328653, 7.325014, 7.328701, 
    7.310239, 7.318144, 7.301918, 7.238967, 7.257422, 7.202482, 7.169594, 
    7.147838, 7.132425, 7.134602, 7.138752, 7.160122, 7.180268, 7.195649, 
    7.205951, 7.216115, 7.246926, 7.263293, 7.300026, 7.293395, 7.304638, 
    7.315402, 7.333492, 7.330513, 7.33849, 7.304347, 7.327022, 7.289618, 
    7.299832, 7.218851, 7.188221, 7.175209, 7.163856, 7.136276, 7.155312, 
    7.147802, 7.165684, 7.177061, 7.171434, 7.206233, 7.192687, 7.264264, 
    7.233366, 7.314146, 7.294756, 7.3188, 7.306525, 7.327566, 7.308627, 
    7.341463, 7.348625, 7.343729, 7.362557, 7.307578, 7.32865, 7.171275, 
    7.172192, 7.17647, 7.157678, 7.156531, 7.139355, 7.154639, 7.161154, 
    7.177723, 7.187534, 7.196871, 7.217436, 7.240454, 7.272744, 7.296011, 
    7.311638, 7.302055, 7.310515, 7.301057, 7.296628, 7.345939, 7.318216, 
    7.359847, 7.35754, 7.338679, 7.3578, 7.172837, 7.167558, 7.149244, 
    7.163573, 7.137487, 7.152075, 7.160473, 7.192964, 7.200125, 7.206761, 
    7.21989, 7.236763, 7.266434, 7.292327, 7.31603, 7.314291, 7.314903, 
    7.320203, 7.307077, 7.32236, 7.324924, 7.318216, 7.357231, 7.346068, 
    7.357491, 7.350222, 7.169274, 7.178162, 7.173357, 7.182392, 7.176024, 
    7.204367, 7.212883, 7.252841, 7.236428, 7.262571, 7.239083, 7.243239, 
    7.263413, 7.240353, 7.290893, 7.256588, 7.320409, 7.286039, 7.322566, 
    7.315927, 7.326925, 7.336782, 7.349204, 7.372157, 7.366838, 7.386071, 
    7.191431, 7.202987, 7.201974, 7.214086, 7.223052, 7.242523, 7.273831, 
    7.262047, 7.283696, 7.288045, 7.255164, 7.275335, 7.210733, 7.221134, 
    7.214944, 7.192339, 7.264754, 7.227516, 7.296395, 7.276142, 7.335375, 
    7.305865, 7.36391, 7.388819, 7.412346, 7.439885, 7.209305, 7.201446, 
    7.215528, 7.235039, 7.253193, 7.277375, 7.279855, 7.284391, 7.296156, 
    7.306057, 7.28582, 7.308541, 7.223538, 7.267995, 7.198472, 7.219344, 
    7.23389, 7.227511, 7.260703, 7.268541, 7.300452, 7.283947, 7.382661, 
    7.338859, 7.460922, 7.426652, 7.1987, 7.209281, 7.246194, 7.228613, 
    7.278994, 7.291431, 7.301558, 7.314512, 7.315916, 7.3236, 7.31101, 
    7.323105, 7.277427, 7.297812, 7.241974, 7.255532, 7.249294, 7.242453, 
    7.263583, 7.286137, 7.286628, 7.293869, 7.314289, 7.279199, 7.388313, 
    7.320763, 7.220832, 7.241262, 7.244194, 7.23627, 7.290183, 7.270614, 
    7.323414, 7.309117, 7.332556, 7.320901, 7.319187, 7.304243, 7.294949, 
    7.271509, 7.252479, 7.237421, 7.24092, 7.257469, 7.28752, 7.316039, 
    7.309783, 7.330773, 7.275332, 7.298535, 7.289558, 7.312986, 7.261733, 
    7.305335, 7.250615, 7.255402, 7.270226, 7.300106, 7.306741, 7.313816, 
    7.309452, 7.288286, 7.284826, 7.269867, 7.265736, 7.25436, 7.244949, 
    7.253545, 7.26258, 7.288298, 7.311527, 7.336921, 7.34315, 7.372906, 
    7.348665, 7.388689, 7.354633, 7.413672, 7.30788, 7.35365, 7.270904, 
    7.279787, 7.295863, 7.332857, 7.312876, 7.336252, 7.284691, 7.258037, 
    7.251163, 7.238334, 7.251456, 7.250389, 7.26296, 7.258919, 7.289153, 
    7.272902, 7.319141, 7.33607, 7.38405, 7.413578, 7.443741, 7.457083, 
    7.461148, 7.462848 ;

 WIND =
  5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932 ;

 WOODC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 WOODC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOODC_LOSS =
  1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11 ;

 WOOD_HARVESTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOOD_HARVESTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WTGQ =
  0.0002557223, 0.0002556714, 0.0002556811, 0.0002556405, 0.0002556627, 
    0.0002556364, 0.0002557116, 0.0002556697, 0.0002556962, 0.0002557172, 
    0.0002555632, 0.0002556386, 0.0002554812, 0.0002555298, 0.0002554067, 
    0.0002554893, 0.00025539, 0.0002554082, 0.0002553511, 0.0002553674, 
    0.0002552963, 0.0002553436, 0.0002552581, 0.0002553071, 0.0002552998, 
    0.0002553453, 0.0002556226, 0.0002555728, 0.0002556257, 0.0002556186, 
    0.0002556216, 0.0002556625, 0.0002556838, 0.0002557256, 0.0002557179, 
    0.0002556868, 0.0002556153, 0.000255639, 0.0002555777, 0.000255579, 
    0.0002555115, 0.000255542, 0.0002554281, 0.0002554602, 0.0002553667, 
    0.0002553903, 0.000255368, 0.0002553746, 0.0002553679, 0.0002554025, 
    0.0002553877, 0.0002554179, 0.0002555364, 0.0002555018, 0.0002556056, 
    0.0002556696, 0.00025571, 0.0002557393, 0.0002557351, 0.0002557274, 
    0.0002556866, 0.0002556476, 0.0002556182, 0.0002555986, 0.0002555792, 
    0.000255523, 0.0002554914, 0.000255422, 0.0002554338, 0.0002554133, 
    0.0002553927, 0.000255359, 0.0002553645, 0.0002553498, 0.0002554133, 
    0.0002553714, 0.0002554407, 0.0002554218, 0.000255577, 0.0002556325, 
    0.0002556587, 0.0002556793, 0.000255732, 0.0002556958, 0.0002557101, 
    0.0002556754, 0.0002556538, 0.0002556643, 0.0002555981, 0.0002556239, 
    0.0002554895, 0.0002555473, 0.000255395, 0.0002554313, 0.0002553863, 
    0.0002554091, 0.0002553702, 0.0002554052, 0.0002553442, 0.0002553313, 
    0.0002553402, 0.0002553049, 0.0002554072, 0.0002553683, 0.0002556648, 
    0.0002556631, 0.0002556548, 0.0002556913, 0.0002556934, 0.000255726, 
    0.0002556967, 0.0002556845, 0.0002556523, 0.0002556338, 0.0002556161, 
    0.000255577, 0.000255534, 0.0002554731, 0.000255429, 0.0002553995, 
    0.0002554174, 0.0002554017, 0.0002554193, 0.0002554275, 0.0002553363, 
    0.0002553877, 0.00025531, 0.0002553142, 0.0002553496, 0.0002553137, 
    0.0002556618, 0.0002556717, 0.0002557071, 0.0002556794, 0.0002557295, 
    0.0002557019, 0.0002556862, 0.0002556241, 0.0002556097, 0.0002555973, 
    0.0002555722, 0.0002555404, 0.0002554849, 0.0002554362, 0.0002553913, 
    0.0002553946, 0.0002553934, 0.0002553837, 0.0002554082, 0.0002553797, 
    0.0002553752, 0.0002553874, 0.0002553148, 0.0002553355, 0.0002553143, 
    0.0002553277, 0.0002556684, 0.0002556516, 0.0002556607, 0.0002556437, 
    0.000255656, 0.0002556026, 0.0002555866, 0.000255511, 0.0002555412, 
    0.0002554923, 0.000255536, 0.0002555284, 0.000255492, 0.0002555334, 
    0.0002554394, 0.0002555043, 0.0002553833, 0.0002554492, 0.0002553793, 
    0.0002553915, 0.000255371, 0.000255353, 0.0002553297, 0.0002552877, 
    0.0002552973, 0.0002552618, 0.0002556263, 0.0002556048, 0.0002556061, 
    0.0002555832, 0.0002555665, 0.0002555294, 0.0002554707, 0.0002554926, 
    0.0002554519, 0.0002554439, 0.0002555055, 0.0002554682, 0.00025559, 
    0.0002555709, 0.0002555818, 0.0002556249, 0.0002554884, 0.0002555587, 
    0.0002554284, 0.0002554663, 0.0002553556, 0.0002554112, 0.0002553028, 
    0.000255258, 0.0002552132, 0.0002551641, 0.0002555925, 0.0002556071, 
    0.0002555804, 0.0002555444, 0.0002555095, 0.0002554641, 0.0002554591, 
    0.0002554508, 0.0002554285, 0.00025541, 0.0002554487, 0.0002554053, 
    0.0002555676, 0.000255482, 0.0002556132, 0.0002555744, 0.0002555463, 
    0.000255558, 0.000255495, 0.0002554803, 0.0002554211, 0.0002554514, 
    0.0002552695, 0.0002553499, 0.0002551248, 0.000255188, 0.0002556124, 
    0.0002555922, 0.0002555231, 0.0002555559, 0.0002554607, 0.0002554376, 
    0.0002554183, 0.0002553946, 0.0002553916, 0.0002553775, 0.0002554007, 
    0.0002553782, 0.000255464, 0.0002554255, 0.0002555303, 0.0002555051, 
    0.0002555165, 0.0002555294, 0.0002554896, 0.0002554482, 0.0002554464, 
    0.0002554333, 0.000255398, 0.0002554603, 0.0002552608, 0.0002553855, 
    0.0002555703, 0.0002555329, 0.0002555264, 0.0002555411, 0.00025544, 
    0.0002554767, 0.0002553777, 0.0002554043, 0.0002553606, 0.0002553824, 
    0.0002553856, 0.0002554134, 0.0002554309, 0.0002554752, 0.0002555109, 
    0.0002555389, 0.0002555323, 0.0002555016, 0.0002554455, 0.0002553918, 
    0.0002554037, 0.0002553639, 0.0002554677, 0.0002554246, 0.0002554415, 
    0.0002553972, 0.0002554934, 0.0002554142, 0.000255514, 0.000255505, 
    0.0002554774, 0.0002554223, 0.0002554087, 0.0002553959, 0.0002554036, 
    0.0002554439, 0.0002554501, 0.0002554778, 0.000255486, 0.0002555069, 
    0.0002555247, 0.0002555087, 0.0002554921, 0.0002554435, 0.0002554003, 
    0.0002553528, 0.0002553409, 0.0002552879, 0.0002553323, 0.0002552603, 
    0.0002553234, 0.0002552133, 0.0002554083, 0.0002553234, 0.0002554758, 
    0.0002554592, 0.00025543, 0.0002553612, 0.0002553974, 0.0002553547, 
    0.0002554502, 0.000255501, 0.000255513, 0.0002555373, 0.0002555125, 
    0.0002555145, 0.0002554907, 0.0002554983, 0.0002554418, 0.0002554721, 
    0.0002553859, 0.0002553548, 0.0002552658, 0.000255212, 0.0002551558, 
    0.0002551314, 0.0002551239, 0.0002551209 ;

 W_SCALAR =
  0.6261148, 0.627772, 0.62745, 0.6287856, 0.6280448, 0.6289191, 0.6264508, 
    0.6278378, 0.6269525, 0.626264, 0.6313739, 0.6288451, 0.6339946, 
    0.6323858, 0.6364231, 0.6337445, 0.6369624, 0.6363456, 0.6382005, 
    0.6376694, 0.6400391, 0.6384455, 0.6412655, 0.6396586, 0.6399102, 
    0.6383929, 0.6293542, 0.6310594, 0.6292531, 0.6294965, 0.6293873, 
    0.6280602, 0.627391, 0.6259879, 0.6262427, 0.6272731, 0.6296058, 
    0.6288143, 0.6308079, 0.6307629, 0.6329789, 0.6319802, 0.6356989, 
    0.6346431, 0.6376916, 0.6369256, 0.6376556, 0.6374343, 0.6376585, 
    0.636535, 0.6370165, 0.6360273, 0.6321673, 0.633303, 0.629913, 0.6278706, 
    0.6265118, 0.6255469, 0.6256833, 0.6259434, 0.6272792, 0.6285336, 
    0.6294889, 0.6301275, 0.6307564, 0.6326588, 0.633664, 0.6359124, 
    0.6355067, 0.6361938, 0.6368494, 0.6379496, 0.6377686, 0.6382532, 
    0.6361755, 0.6375567, 0.6352757, 0.6359, 0.630928, 0.6290279, 0.62822, 
    0.6275119, 0.6257882, 0.6269789, 0.6265096, 0.6276255, 0.6283342, 
    0.6279837, 0.630145, 0.6293051, 0.6337236, 0.6318223, 0.6367729, 0.63559, 
    0.6370563, 0.6363083, 0.6375897, 0.6364365, 0.6384333, 0.6388679, 
    0.638571, 0.6397107, 0.6363725, 0.6376557, 0.6279739, 0.6280311, 
    0.6282973, 0.6271266, 0.6270549, 0.625981, 0.6269366, 0.6273434, 
    0.6283752, 0.6289852, 0.6295649, 0.6308383, 0.6322592, 0.6342434, 
    0.6356667, 0.63662, 0.6360355, 0.6365516, 0.6359747, 0.6357042, 
    0.6387051, 0.637021, 0.6395468, 0.6394072, 0.6382647, 0.6394229, 
    0.6280712, 0.6277422, 0.6265996, 0.6274939, 0.625864, 0.6267766, 
    0.6273012, 0.6293229, 0.6297665, 0.6301779, 0.6309899, 0.6320313, 
    0.6338563, 0.6354419, 0.6368875, 0.6367816, 0.6368189, 0.6371417, 
    0.636342, 0.6372729, 0.6374292, 0.6370207, 0.6393885, 0.6387125, 
    0.6394042, 0.6389641, 0.6278492, 0.6284026, 0.6281036, 0.6286659, 
    0.6282698, 0.6300302, 0.6305575, 0.6330219, 0.6320109, 0.6336194, 
    0.6321743, 0.6324306, 0.6336721, 0.6322524, 0.6353546, 0.6332525, 
    0.6371542, 0.6350583, 0.6372855, 0.6368812, 0.6375504, 0.6381494, 
    0.6389025, 0.640291, 0.6399696, 0.6411298, 0.6292272, 0.6299443, 
    0.629881, 0.630631, 0.6311855, 0.6323861, 0.6343096, 0.6335866, 
    0.6349136, 0.6351798, 0.6331637, 0.6344021, 0.6304239, 0.6310676, 
    0.6306843, 0.6292838, 0.6337535, 0.6314616, 0.6356903, 0.6344512, 
    0.6380641, 0.6362687, 0.6397927, 0.6412964, 0.6427092, 0.6443588, 
    0.6303353, 0.6298483, 0.6307201, 0.6319257, 0.6330429, 0.6345268, 
    0.6346784, 0.6349562, 0.6356754, 0.6362798, 0.6350442, 0.6364312, 
    0.6312171, 0.6339521, 0.6296642, 0.6309571, 0.6318546, 0.6314608, 
    0.6335039, 0.633985, 0.6359382, 0.6349289, 0.6409255, 0.6382761, 
    0.6456128, 0.6435673, 0.6296781, 0.6303336, 0.6326126, 0.6315288, 
    0.6346257, 0.6353869, 0.6360052, 0.6367954, 0.6368806, 0.6373485, 
    0.6365817, 0.6373182, 0.6345299, 0.6357767, 0.6323522, 0.6331866, 
    0.6328028, 0.6323817, 0.6336808, 0.6350636, 0.635093, 0.6355361, 
    0.6367843, 0.6346382, 0.6412675, 0.6371781, 0.631048, 0.6323094, 
    0.6324891, 0.6320008, 0.6353106, 0.6341124, 0.6373371, 0.6364663, 
    0.6378927, 0.6371841, 0.6370798, 0.6361691, 0.6356018, 0.6341674, 
    0.632999, 0.6320716, 0.6322873, 0.6333058, 0.6351482, 0.6368884, 
    0.6365075, 0.6377843, 0.6344014, 0.6358212, 0.6352727, 0.6367022, 
    0.6335675, 0.6362381, 0.632884, 0.6331784, 0.6340886, 0.6359175, 
    0.6363215, 0.6367531, 0.6364867, 0.6351948, 0.634983, 0.6340664, 
    0.6338133, 0.6331143, 0.6325353, 0.6330644, 0.6336197, 0.6351953, 
    0.6366136, 0.638158, 0.6385356, 0.6403375, 0.6388711, 0.6412902, 
    0.6392343, 0.6427908, 0.6363924, 0.6391734, 0.6341299, 0.6346742, 
    0.6356583, 0.6379119, 0.6366956, 0.6381178, 0.6349747, 0.633341, 
    0.6329178, 0.6321281, 0.6329358, 0.6328701, 0.6336426, 0.6333944, 
    0.6352476, 0.6342525, 0.6370773, 0.6381066, 0.6410084, 0.6427839, 
    0.6445881, 0.6453838, 0.6456259, 0.6457272,
  0.5467909, 0.548835, 0.5484377, 0.5500853, 0.5491714, 0.5502501, 0.5472054, 
    0.5489162, 0.5478241, 0.5469749, 0.5532789, 0.5501587, 0.5565134, 
    0.5545277, 0.5595115, 0.5562047, 0.5601775, 0.5594159, 0.5617064, 
    0.5610505, 0.5639775, 0.5620091, 0.5654924, 0.5635074, 0.5638182, 
    0.5619441, 0.5507868, 0.5528908, 0.5506622, 0.5509623, 0.5508276, 
    0.5491904, 0.5483649, 0.5466344, 0.5469487, 0.5482196, 0.5510973, 
    0.5501208, 0.5525804, 0.5525249, 0.5552596, 0.5540271, 0.5586174, 
    0.5573139, 0.5610779, 0.5601321, 0.5610335, 0.5607602, 0.5610371, 
    0.5596497, 0.5602443, 0.5590229, 0.554258, 0.5556598, 0.5514762, 
    0.5489565, 0.5472805, 0.5460905, 0.5462587, 0.5465795, 0.548227, 
    0.5497745, 0.550953, 0.5517409, 0.5525169, 0.5548645, 0.5561053, 
    0.558881, 0.5583802, 0.5592284, 0.560038, 0.5613967, 0.5611731, 
    0.5617715, 0.5592058, 0.5609115, 0.5580949, 0.5588657, 0.5527286, 
    0.5503842, 0.5493875, 0.5485141, 0.5463881, 0.5478566, 0.5472779, 
    0.5486543, 0.5495284, 0.549096, 0.5517624, 0.5507263, 0.5561789, 
    0.5538322, 0.5599436, 0.558483, 0.5602934, 0.5593698, 0.5609521, 
    0.5595281, 0.5619941, 0.5625306, 0.562164, 0.5635718, 0.5594491, 
    0.5610336, 0.549084, 0.5491545, 0.5494829, 0.5480388, 0.5479504, 
    0.5466259, 0.5478045, 0.5483062, 0.549579, 0.5503316, 0.5510467, 
    0.552618, 0.5543715, 0.5568205, 0.5585777, 0.5597547, 0.559033, 
    0.5596702, 0.5589579, 0.558624, 0.5623296, 0.5602499, 0.5633693, 
    0.5631968, 0.5617857, 0.5632163, 0.549204, 0.5487982, 0.5473888, 
    0.5484918, 0.5464815, 0.5476072, 0.5482541, 0.5507481, 0.5512955, 
    0.5518031, 0.552805, 0.5540902, 0.5563427, 0.5583001, 0.560085, 
    0.5599543, 0.5600003, 0.5603989, 0.5594115, 0.5605609, 0.5607539, 
    0.5602496, 0.5631738, 0.5623388, 0.5631932, 0.5626496, 0.5489301, 
    0.5496128, 0.5492439, 0.5499375, 0.549449, 0.5516208, 0.5522714, 
    0.5553128, 0.554065, 0.5560502, 0.5542667, 0.5545829, 0.5561153, 
    0.5543631, 0.5581924, 0.5555974, 0.5604144, 0.5578266, 0.5605764, 
    0.5600773, 0.5609036, 0.5616434, 0.5625735, 0.5642887, 0.5638916, 
    0.5653248, 0.5506301, 0.5515149, 0.5514368, 0.5523622, 0.5530463, 
    0.5545281, 0.5569023, 0.5560098, 0.5576478, 0.5579765, 0.5554878, 
    0.5570164, 0.5521066, 0.5529009, 0.5524279, 0.5506999, 0.5562158, 
    0.5533872, 0.5586067, 0.5570769, 0.561538, 0.559321, 0.563673, 0.5655306, 
    0.5672763, 0.5693149, 0.5519974, 0.5513964, 0.5524722, 0.5539598, 
    0.5553386, 0.5571703, 0.5573575, 0.5577005, 0.5585884, 0.5593346, 
    0.5578091, 0.5595216, 0.5530853, 0.556461, 0.5511693, 0.5527645, 
    0.5538721, 0.5533862, 0.5559078, 0.5565016, 0.5589129, 0.5576667, 
    0.5650725, 0.5617998, 0.5708649, 0.5683366, 0.5511864, 0.5519952, 
    0.5548077, 0.55347, 0.5572925, 0.5582322, 0.5589957, 0.5599713, 
    0.5600765, 0.5606543, 0.5597074, 0.5606169, 0.5571742, 0.5587134, 
    0.5544862, 0.5555161, 0.5550423, 0.5545226, 0.5561261, 0.5578331, 
    0.5578694, 0.5584164, 0.5599575, 0.5573079, 0.5654948, 0.5604437, 
    0.5528768, 0.5544333, 0.5546553, 0.5540525, 0.558138, 0.5566588, 
    0.5606402, 0.5595649, 0.5613263, 0.5604513, 0.5603225, 0.559198, 
    0.5584975, 0.5567267, 0.5552845, 0.55414, 0.5544061, 0.5556632, 
    0.5579374, 0.5600861, 0.5596157, 0.5611925, 0.5570156, 0.5587683, 
    0.5580912, 0.5598563, 0.5559862, 0.5592831, 0.5551426, 0.5555059, 
    0.5566294, 0.5588874, 0.5593861, 0.559919, 0.5595902, 0.5579951, 
    0.5577335, 0.5566021, 0.5562897, 0.5554268, 0.5547122, 0.5553652, 
    0.5560507, 0.5579957, 0.5597468, 0.561654, 0.5621203, 0.564346, 
    0.5625347, 0.565523, 0.5629832, 0.567377, 0.5594736, 0.562908, 0.5566804, 
    0.5573523, 0.5585672, 0.56135, 0.559848, 0.5616044, 0.5577233, 0.5557066, 
    0.5551842, 0.5542096, 0.5552065, 0.5551254, 0.5560789, 0.5557725, 
    0.5580602, 0.5568317, 0.5603194, 0.5615904, 0.5651748, 0.5673686, 
    0.5695983, 0.5705819, 0.5708812, 0.5710062,
  0.5141823, 0.5164323, 0.515995, 0.5178089, 0.5168027, 0.5179903, 0.5146385, 
    0.5165216, 0.5153195, 0.5143847, 0.521326, 0.5178897, 0.52489, 0.5227019, 
    0.5281949, 0.5245497, 0.5289292, 0.5280896, 0.5306154, 0.529892, 
    0.5331206, 0.5309492, 0.5347923, 0.5326021, 0.532945, 0.5308776, 
    0.5185813, 0.5208985, 0.5184441, 0.5187746, 0.5186262, 0.5168235, 
    0.5159149, 0.5140101, 0.514356, 0.5157548, 0.5189232, 0.5178479, 
    0.5205567, 0.5204955, 0.5235084, 0.5221503, 0.5272092, 0.5257723, 
    0.5299222, 0.5288792, 0.5298733, 0.5295719, 0.5298772, 0.5283473, 
    0.5290029, 0.5276563, 0.5224048, 0.5239493, 0.5193405, 0.516566, 
    0.5147212, 0.5134115, 0.5135967, 0.5139497, 0.515763, 0.5174666, 
    0.5187643, 0.519632, 0.5204868, 0.523073, 0.5244403, 0.5274998, 
    0.5269477, 0.5278828, 0.5287754, 0.5302737, 0.5300272, 0.5306872, 
    0.5278579, 0.5297386, 0.5266332, 0.5274829, 0.5207199, 0.518138, 
    0.5170406, 0.5160791, 0.513739, 0.5153552, 0.5147182, 0.5162333, 
    0.5171957, 0.5167197, 0.5196558, 0.5185147, 0.5245213, 0.5219356, 
    0.5286713, 0.527061, 0.5290571, 0.5280387, 0.5297835, 0.5282132, 
    0.5309327, 0.5315245, 0.5311201, 0.5326731, 0.5281262, 0.5298734, 
    0.5167064, 0.5167841, 0.5171456, 0.5155559, 0.5154586, 0.5140007, 
    0.5152978, 0.5158501, 0.5172514, 0.5180801, 0.5188676, 0.5205981, 
    0.5225298, 0.5252284, 0.5271654, 0.5284631, 0.5276674, 0.5283699, 
    0.5275846, 0.5272164, 0.5313028, 0.5290091, 0.5324497, 0.5322595, 
    0.5307029, 0.5322809, 0.5168386, 0.5163918, 0.5148403, 0.5160546, 
    0.5138418, 0.5150807, 0.5157929, 0.5185387, 0.5191414, 0.5197005, 
    0.5208041, 0.5222199, 0.5247018, 0.5268593, 0.5288273, 0.5286831, 
    0.5287339, 0.5291734, 0.5280847, 0.5293521, 0.5295649, 0.5290087, 
    0.532234, 0.5313129, 0.5322554, 0.5316557, 0.516537, 0.5172886, 
    0.5168825, 0.5176462, 0.5171083, 0.5194997, 0.5202163, 0.5235668, 
    0.5221921, 0.5243795, 0.5224143, 0.5227627, 0.5244512, 0.5225205, 
    0.5267406, 0.5238805, 0.5291905, 0.5263373, 0.5293692, 0.5288188, 
    0.52973, 0.5305459, 0.5315718, 0.533464, 0.5330259, 0.5346074, 0.5184087, 
    0.5193831, 0.5192971, 0.5203164, 0.5210699, 0.5227023, 0.5253186, 
    0.524335, 0.5261403, 0.5265027, 0.5237598, 0.5254443, 0.5200348, 
    0.5209097, 0.5203887, 0.5184857, 0.5245619, 0.5214453, 0.5271974, 
    0.5255111, 0.5304296, 0.5279849, 0.5327848, 0.5348344, 0.5367613, 
    0.539012, 0.5199145, 0.5192527, 0.5204375, 0.5220762, 0.5235954, 
    0.525614, 0.5258204, 0.5261984, 0.5271772, 0.5279999, 0.5263181, 
    0.5282061, 0.5211129, 0.5248322, 0.5190026, 0.5207595, 0.5219796, 
    0.5214443, 0.5242226, 0.524877, 0.527535, 0.5261612, 0.5343289, 
    0.5307184, 0.5407239, 0.5379319, 0.5190214, 0.5199122, 0.5230103, 
    0.5215366, 0.5257487, 0.5267845, 0.5276262, 0.5287019, 0.5288179, 
    0.5294551, 0.5284109, 0.5294138, 0.5256183, 0.5273151, 0.5226561, 
    0.523791, 0.5232689, 0.5226963, 0.5244632, 0.5263446, 0.5263845, 
    0.5269876, 0.5286866, 0.5257657, 0.534795, 0.5292228, 0.5208831, 
    0.5225978, 0.5228423, 0.5221784, 0.5266807, 0.5250502, 0.5294395, 
    0.5282539, 0.5301961, 0.5292312, 0.5290892, 0.5278493, 0.527077, 
    0.5251251, 0.5235357, 0.5222747, 0.5225679, 0.523953, 0.5264596, 
    0.5288286, 0.5283098, 0.5300485, 0.5254434, 0.5273756, 0.526629, 
    0.5285751, 0.5243089, 0.527943, 0.5233794, 0.5237797, 0.5250179, 
    0.5275068, 0.5280567, 0.5286442, 0.5282816, 0.5265232, 0.5262348, 
    0.5249877, 0.5246434, 0.5236925, 0.5229052, 0.5236247, 0.52438, 
    0.5265238, 0.5284544, 0.5305575, 0.5310718, 0.5335273, 0.531529, 
    0.534826, 0.5320237, 0.5368724, 0.5281531, 0.5319408, 0.5250741, 
    0.5258147, 0.5271538, 0.5302223, 0.5285659, 0.5305029, 0.5262235, 
    0.5240009, 0.5234252, 0.5223514, 0.5234498, 0.5233604, 0.5244111, 
    0.5240735, 0.5265949, 0.5252408, 0.5290857, 0.5304875, 0.5344418, 
    0.5368631, 0.539325, 0.5404113, 0.5407418, 0.54088,
  0.507082, 0.5094726, 0.5090079, 0.5109358, 0.5098663, 0.5111287, 0.5075666, 
    0.5095676, 0.5082902, 0.5072972, 0.5146762, 0.5110217, 0.5184694, 
    0.5161402, 0.5219896, 0.5181071, 0.5227723, 0.5218774, 0.5245696, 
    0.5237985, 0.5272414, 0.5249255, 0.5290251, 0.5266883, 0.527054, 
    0.5248492, 0.5117571, 0.5142214, 0.5116111, 0.5119625, 0.5118048, 
    0.5098885, 0.5089228, 0.5068991, 0.5072665, 0.5087527, 0.5121205, 
    0.5109773, 0.5138578, 0.5137928, 0.5169986, 0.5155533, 0.5209395, 
    0.5194089, 0.5238306, 0.5227189, 0.5237784, 0.5234572, 0.5237826, 
    0.5221521, 0.5228508, 0.5214157, 0.515824, 0.5174679, 0.5125643, 
    0.5096148, 0.5076545, 0.5062633, 0.50646, 0.506835, 0.5087614, 0.510572, 
    0.5119516, 0.5128743, 0.5137834, 0.5165351, 0.5179906, 0.521249, 
    0.5206609, 0.521657, 0.5226083, 0.5242054, 0.5239425, 0.5246461, 
    0.5216306, 0.5236349, 0.5203258, 0.5212311, 0.5140314, 0.5112857, 
    0.5101191, 0.5090972, 0.5066112, 0.5083281, 0.5076514, 0.5092612, 
    0.510284, 0.5097781, 0.5128996, 0.5116862, 0.5180768, 0.5153248, 
    0.5224974, 0.5207816, 0.5229085, 0.5218232, 0.5236828, 0.5220092, 
    0.5249079, 0.525539, 0.5251077, 0.526764, 0.5219164, 0.5237786, 0.509764, 
    0.5098465, 0.5102308, 0.5085413, 0.5084379, 0.5068891, 0.5082672, 
    0.508854, 0.5103432, 0.5112241, 0.5120614, 0.5139019, 0.5159571, 
    0.5188298, 0.5208928, 0.5222754, 0.5214276, 0.5221761, 0.5213394, 
    0.5209472, 0.5253026, 0.5228573, 0.5265257, 0.5263228, 0.5246629, 
    0.5263457, 0.5099044, 0.5094296, 0.5077811, 0.5090712, 0.5067204, 
    0.5080364, 0.5087932, 0.5117117, 0.5123526, 0.5129471, 0.514121, 
    0.5156273, 0.5182691, 0.5205668, 0.5226636, 0.5225099, 0.5225641, 
    0.5230325, 0.5218722, 0.5232229, 0.5234497, 0.522857, 0.5262956, 
    0.5253134, 0.5263185, 0.5256789, 0.5095839, 0.5103828, 0.5099511, 
    0.5107629, 0.5101911, 0.5127336, 0.5134957, 0.5170608, 0.5155977, 
    0.5179259, 0.5158342, 0.5162049, 0.5180022, 0.5159472, 0.5204403, 
    0.5173947, 0.5230507, 0.5200107, 0.5232412, 0.5226545, 0.5236257, 
    0.5244955, 0.5255894, 0.5276077, 0.5271404, 0.5288278, 0.5115736, 
    0.5126095, 0.5125182, 0.5136021, 0.5144038, 0.5161406, 0.5189258, 
    0.5178785, 0.5198009, 0.5201868, 0.5172662, 0.5190597, 0.5133027, 
    0.5142333, 0.5136791, 0.5116554, 0.5181201, 0.5148032, 0.520927, 
    0.5191308, 0.5243715, 0.5217658, 0.5268831, 0.5290701, 0.531127, 
    0.5335308, 0.5131748, 0.5124709, 0.513731, 0.5154744, 0.5170912, 
    0.5192404, 0.5194601, 0.5198628, 0.5209053, 0.5217819, 0.5199902, 
    0.5220016, 0.5144494, 0.5184079, 0.5122049, 0.5140735, 0.5153716, 
    0.514802, 0.5177588, 0.5184556, 0.5212865, 0.5198231, 0.5285305, 
    0.5246794, 0.5353601, 0.532377, 0.512225, 0.5131723, 0.5164685, 
    0.5149003, 0.5193838, 0.5204871, 0.5213837, 0.52253, 0.5226536, 
    0.5233327, 0.5222199, 0.5232886, 0.519245, 0.5210522, 0.5160915, 
    0.5172994, 0.5167437, 0.5161343, 0.518015, 0.5200185, 0.520061, 
    0.5207034, 0.5225136, 0.5194019, 0.5290279, 0.5230851, 0.5142051, 
    0.5160295, 0.5162897, 0.5155831, 0.5203764, 0.51864, 0.523316, 0.5220525, 
    0.5241226, 0.5230941, 0.5229427, 0.5216213, 0.5207987, 0.5187197, 
    0.5170277, 0.5156856, 0.5159976, 0.5174718, 0.5201409, 0.5226649, 
    0.5221121, 0.5239653, 0.5190588, 0.5211167, 0.5203214, 0.5223948, 
    0.5178508, 0.5217212, 0.5168613, 0.5172874, 0.5186055, 0.5212564, 
    0.5218424, 0.5224685, 0.5220821, 0.5202087, 0.5199016, 0.5185735, 
    0.5182068, 0.5171946, 0.5163566, 0.5171223, 0.5179265, 0.5202093, 
    0.5222661, 0.5245079, 0.5250563, 0.5276752, 0.5255437, 0.5290611, 
    0.5260714, 0.5312456, 0.5219451, 0.5259829, 0.5186654, 0.5194541, 
    0.5208805, 0.5241506, 0.5223851, 0.5244496, 0.5198895, 0.5175229, 
    0.5169101, 0.5157672, 0.5169362, 0.5168411, 0.5179596, 0.5176002, 
    0.5202851, 0.518843, 0.522939, 0.5244332, 0.5286511, 0.5312357, 
    0.5338653, 0.535026, 0.5353792, 0.5355269,
  0.5310288, 0.5334982, 0.5330179, 0.5350106, 0.533905, 0.5352101, 0.5315292, 
    0.5335963, 0.5322765, 0.5312509, 0.5388809, 0.5350995, 0.5428115, 
    0.5403972, 0.5464646, 0.5424359, 0.5472774, 0.546348, 0.5491452, 
    0.5483436, 0.5519241, 0.5495152, 0.5537811, 0.5513485, 0.5517291, 
    0.5494357, 0.5358599, 0.53841, 0.535709, 0.5360725, 0.5359093, 0.5339279, 
    0.53293, 0.5308399, 0.5312192, 0.5327542, 0.5362359, 0.5350536, 
    0.5380336, 0.5379663, 0.5412867, 0.5397893, 0.5453742, 0.543786, 
    0.548377, 0.547222, 0.5483229, 0.547989, 0.5483272, 0.5466332, 0.5473589, 
    0.5458686, 0.5400698, 0.5417732, 0.536695, 0.533645, 0.5316199, 
    0.5301836, 0.5303866, 0.5307737, 0.5327632, 0.5346345, 0.5360612, 
    0.5370158, 0.5379566, 0.5408065, 0.5423151, 0.5456956, 0.5450851, 
    0.5461192, 0.5471071, 0.5487666, 0.5484933, 0.5492247, 0.5460917, 
    0.5481737, 0.5447374, 0.545677, 0.5382133, 0.5353725, 0.5341663, 
    0.5331103, 0.5305427, 0.5323157, 0.5316167, 0.5332797, 0.5343368, 
    0.5338139, 0.5370419, 0.5357866, 0.5424045, 0.5395526, 0.5469918, 
    0.5452104, 0.547419, 0.5462918, 0.5482234, 0.5464849, 0.5494968, 
    0.5501531, 0.5497046, 0.5514273, 0.5463886, 0.5483229, 0.5337992, 
    0.5338845, 0.5342818, 0.5325359, 0.5324291, 0.5308296, 0.5322527, 
    0.532859, 0.534398, 0.5353088, 0.5361747, 0.5380793, 0.5402075, 
    0.5431852, 0.5453258, 0.5467614, 0.545881, 0.5466582, 0.5457894, 
    0.5453822, 0.5499072, 0.5473658, 0.5511795, 0.5509683, 0.5492421, 
    0.5509921, 0.5339444, 0.5334537, 0.5317506, 0.5330834, 0.5306554, 
    0.5320144, 0.5327961, 0.5358131, 0.536476, 0.5370911, 0.5383061, 
    0.5398659, 0.5426038, 0.5449874, 0.5471645, 0.5470049, 0.5470611, 
    0.5475478, 0.5463426, 0.5477456, 0.5479812, 0.5473654, 0.55094, 
    0.5499184, 0.5509638, 0.5502986, 0.5336131, 0.5344389, 0.5339927, 
    0.5348319, 0.5342407, 0.5368702, 0.5376589, 0.5413513, 0.5398353, 
    0.542248, 0.5400802, 0.5404643, 0.5423271, 0.5401973, 0.5448561, 
    0.5416973, 0.5475667, 0.5444103, 0.5477645, 0.5471551, 0.5481641, 
    0.5490681, 0.5502055, 0.5523053, 0.551819, 0.5535756, 0.5356702, 
    0.5367419, 0.5366473, 0.537769, 0.5385988, 0.5403978, 0.5432849, 
    0.5421989, 0.5441927, 0.5445932, 0.5415641, 0.5434238, 0.5374591, 
    0.5384223, 0.5378487, 0.5357548, 0.5424494, 0.5390124, 0.5453612, 
    0.5434975, 0.5489392, 0.5462322, 0.5515513, 0.5538279, 0.555971, 
    0.5584781, 0.5373267, 0.5365984, 0.5379024, 0.5397075, 0.5413827, 
    0.5436112, 0.5438392, 0.5442569, 0.5453388, 0.5462488, 0.5443891, 
    0.546477, 0.5386461, 0.5427478, 0.5363232, 0.5382569, 0.539601, 
    0.5390112, 0.5420747, 0.5427972, 0.5457345, 0.5442157, 0.553266, 
    0.5492593, 0.5603875, 0.5572744, 0.536344, 0.5373241, 0.5407374, 
    0.5391129, 0.5437599, 0.5449046, 0.5458354, 0.5470257, 0.5471541, 
    0.5478596, 0.5467037, 0.5478138, 0.5436159, 0.5454913, 0.5403469, 
    0.5415985, 0.5410226, 0.5403911, 0.5423404, 0.5444184, 0.5444626, 
    0.5451292, 0.5470088, 0.5437787, 0.553784, 0.5476024, 0.5383931, 
    0.5402825, 0.5405522, 0.5398202, 0.5447899, 0.5429885, 0.5478423, 
    0.5465299, 0.5486805, 0.5476117, 0.5474545, 0.5460821, 0.5452281, 
    0.5430712, 0.5413169, 0.5399263, 0.5402496, 0.5417773, 0.5445455, 
    0.5471659, 0.5465918, 0.548517, 0.5434228, 0.5455582, 0.5447328, 
    0.5468853, 0.5421701, 0.5461859, 0.5411444, 0.5415861, 0.5429527, 
    0.5457033, 0.5463117, 0.5469618, 0.5465606, 0.5446157, 0.5442971, 
    0.5429195, 0.5425393, 0.54149, 0.5406215, 0.541415, 0.5422486, 0.5446165, 
    0.5467517, 0.549081, 0.5496511, 0.5523756, 0.550158, 0.5538185, 
    0.5507067, 0.5560948, 0.5464183, 0.5506147, 0.5430148, 0.5438328, 
    0.545313, 0.5487095, 0.5468752, 0.5490204, 0.5442846, 0.5418302, 
    0.541195, 0.5400109, 0.5412221, 0.5411236, 0.5422829, 0.5419103, 
    0.5446951, 0.543199, 0.5474506, 0.5490034, 0.5533916, 0.5560843, 
    0.558827, 0.5600387, 0.5604075, 0.5605618,
  0.535215, 0.5380583, 0.537505, 0.5398022, 0.5385273, 0.5400323, 0.5357908, 
    0.5381714, 0.5366511, 0.5354705, 0.5442734, 0.5399048, 0.5488272, 
    0.5460286, 0.5530714, 0.5483914, 0.5540173, 0.5529358, 0.5561932, 
    0.555259, 0.5594366, 0.5566247, 0.5616078, 0.5587642, 0.5592087, 
    0.5565321, 0.5407823, 0.5437287, 0.5406081, 0.5410277, 0.5408393, 
    0.5385537, 0.5374036, 0.5349978, 0.5354341, 0.5372012, 0.5412164, 
    0.5398518, 0.5432935, 0.5432156, 0.5470591, 0.5453246, 0.5518034, 
    0.5499582, 0.555298, 0.5539528, 0.5552348, 0.5548459, 0.5552399, 
    0.5532677, 0.5541123, 0.5523782, 0.5456493, 0.5476229, 0.5417466, 
    0.5382276, 0.5358952, 0.5342429, 0.5344764, 0.5349216, 0.5372116, 
    0.5393683, 0.5410146, 0.5421172, 0.5432045, 0.5465026, 0.5482513, 
    0.552177, 0.5514672, 0.5526696, 0.5538191, 0.5557519, 0.5554335, 
    0.5562859, 0.5526377, 0.5550611, 0.5510632, 0.5521553, 0.5435013, 
    0.5402197, 0.5388285, 0.5376113, 0.5346559, 0.5366962, 0.5358915, 
    0.5378065, 0.539025, 0.5384222, 0.5421473, 0.5406978, 0.548355, 
    0.5450506, 0.5536849, 0.5516129, 0.5541821, 0.5528703, 0.555119, 
    0.553095, 0.5566033, 0.5573688, 0.5568456, 0.5588562, 0.5529829, 
    0.555235, 0.5384053, 0.5385036, 0.5389616, 0.5369498, 0.5368267, 
    0.5349858, 0.5366237, 0.5373218, 0.5390956, 0.5401462, 0.5411457, 
    0.5433463, 0.5458089, 0.5492609, 0.5517471, 0.5534167, 0.5523925, 
    0.5532967, 0.5522861, 0.5518126, 0.5570819, 0.5541202, 0.5585667, 
    0.5583202, 0.5563062, 0.558348, 0.5385727, 0.538007, 0.5360457, 
    0.5375804, 0.5347855, 0.5363493, 0.5372494, 0.5407283, 0.5414937, 
    0.5422042, 0.5436085, 0.5454133, 0.5485862, 0.5513538, 0.5538859, 
    0.5537002, 0.5537656, 0.5543321, 0.5529295, 0.5545625, 0.5548369, 
    0.5541198, 0.5582872, 0.557095, 0.558315, 0.5575385, 0.5381908, 
    0.5391428, 0.5386283, 0.539596, 0.5389143, 0.5419489, 0.5428603, 
    0.5471339, 0.5453779, 0.5481735, 0.5456614, 0.5461062, 0.5482653, 
    0.545797, 0.5512012, 0.5475349, 0.5543541, 0.5506833, 0.5545846, 
    0.553875, 0.55505, 0.5561034, 0.55743, 0.559882, 0.5593137, 0.5613673, 
    0.5405633, 0.5418007, 0.5416915, 0.5429876, 0.5439471, 0.5460292, 
    0.5493765, 0.5481166, 0.5504305, 0.5508956, 0.5473805, 0.5495377, 
    0.5426294, 0.543743, 0.5430797, 0.540661, 0.5484071, 0.5444255, 
    0.5517883, 0.5496233, 0.5559531, 0.552801, 0.559001, 0.5616626, 
    0.5641724, 0.5671141, 0.5424764, 0.541635, 0.5431418, 0.54523, 0.5471703, 
    0.5497553, 0.5500199, 0.550505, 0.5517622, 0.5528204, 0.5506586, 
    0.5530857, 0.5440018, 0.5487532, 0.5413172, 0.5435517, 0.5451067, 
    0.5444241, 0.5479726, 0.5488106, 0.5522222, 0.5504572, 0.5610052, 
    0.5563263, 0.5693585, 0.5657009, 0.5413412, 0.5424734, 0.5464225, 
    0.5445418, 0.5499279, 0.5512576, 0.5523396, 0.5537243, 0.5538738, 
    0.5546952, 0.5533496, 0.554642, 0.5497608, 0.5519395, 0.5459703, 
    0.5474204, 0.546753, 0.5460215, 0.5482807, 0.5506927, 0.5507439, 
    0.5515186, 0.5537046, 0.5499498, 0.5616112, 0.5543957, 0.5437092, 
    0.5458958, 0.546208, 0.5453604, 0.5511243, 0.5490325, 0.5546752, 
    0.5531473, 0.5556517, 0.5544065, 0.5542235, 0.5526266, 0.5516335, 
    0.5491284, 0.547094, 0.5454832, 0.5458576, 0.5476277, 0.5508403, 
    0.5538875, 0.5532194, 0.5554611, 0.5495365, 0.5520173, 0.5510579, 
    0.553561, 0.5480832, 0.5527471, 0.5468942, 0.5474061, 0.548991, 0.552186, 
    0.5528935, 0.5536501, 0.5531831, 0.5509219, 0.5505518, 0.5489524, 
    0.5485114, 0.5472946, 0.5462883, 0.5472078, 0.5481742, 0.5509228, 
    0.5534055, 0.5561185, 0.5567833, 0.5599641, 0.5573745, 0.5616516, 
    0.5580149, 0.5643175, 0.5530175, 0.5579075, 0.5490631, 0.5500126, 
    0.5517322, 0.5556855, 0.5535492, 0.5560478, 0.5505372, 0.547689, 
    0.5469528, 0.5455812, 0.5469842, 0.54687, 0.548214, 0.5477819, 0.5510141, 
    0.5492768, 0.554219, 0.5560279, 0.561152, 0.5643053, 0.567524, 0.5689483, 
    0.5693821, 0.5695636,
  0.5840928, 0.5875039, 0.586839, 0.5896026, 0.5880677, 0.5898799, 0.5847825, 
    0.5876399, 0.585814, 0.5843988, 0.5950066, 0.5897262, 0.6005461, 
    0.5971375, 0.6057424, 0.6000144, 0.606905, 0.6055759, 0.6095858, 
    0.6084337, 0.6135982, 0.6101183, 0.6162958, 0.6127648, 0.6133156, 
    0.610004, 0.5907843, 0.5943465, 0.5905741, 0.5910804, 0.5908531, 
    0.5880995, 0.5867173, 0.5838327, 0.5843552, 0.5864743, 0.5913082, 
    0.5896623, 0.5938194, 0.5937251, 0.598391, 0.5962822, 0.6041865, 
    0.6019276, 0.6084818, 0.6068256, 0.6084039, 0.6079248, 0.6084102, 
    0.6059834, 0.6070218, 0.6048915, 0.5966766, 0.5990776, 0.5919484, 
    0.5877073, 0.5849076, 0.5829297, 0.5832089, 0.5837415, 0.5864867, 
    0.58908, 0.5910646, 0.5923963, 0.5937116, 0.5977138, 0.5998436, 
    0.6046446, 0.6037745, 0.605249, 0.6066612, 0.6090413, 0.6086487, 
    0.6097001, 0.6052099, 0.6081898, 0.6032797, 0.6046181, 0.594071, 
    0.5901058, 0.5884302, 0.5869668, 0.5834237, 0.5858681, 0.5849032, 
    0.5872012, 0.5886666, 0.5879413, 0.5924328, 0.5906823, 0.59997, 
    0.5959496, 0.6064963, 0.603953, 0.6071077, 0.6054955, 0.6082612, 
    0.6057714, 0.6100919, 0.6110377, 0.6103912, 0.6128787, 0.6056337, 
    0.608404, 0.5879211, 0.5880393, 0.5885903, 0.5861724, 0.5860248, 
    0.5838185, 0.5857811, 0.5866191, 0.5887516, 0.5900171, 0.5912229, 
    0.5938833, 0.5968704, 0.6010756, 0.6041175, 0.6061666, 0.6049091, 
    0.6060191, 0.6047784, 0.6041979, 0.6106832, 0.6070316, 0.6125202, 
    0.6122149, 0.6097252, 0.6122493, 0.5881223, 0.5874423, 0.585088, 
    0.5869296, 0.5835787, 0.585452, 0.5865321, 0.590719, 0.591643, 0.5925015, 
    0.5942009, 0.5963899, 0.600252, 0.6036355, 0.6067434, 0.606515, 
    0.6065955, 0.6072922, 0.6055682, 0.6075758, 0.6079137, 0.607031, 
    0.612174, 0.6106994, 0.6122084, 0.6112477, 0.5876632, 0.5888084, 
    0.5881893, 0.5893542, 0.5885333, 0.592193, 0.593295, 0.598482, 0.5963469, 
    0.5997487, 0.5966913, 0.5972319, 0.5998606, 0.596856, 0.6034486, 
    0.5989705, 0.6073194, 0.6028146, 0.607603, 0.6067299, 0.6081761, 
    0.6094749, 0.6111134, 0.614151, 0.6134459, 0.6159967, 0.59052, 0.5920138, 
    0.5918819, 0.5934491, 0.5946111, 0.5971382, 0.6012169, 0.5996793, 
    0.6025052, 0.6030745, 0.5987824, 0.6014137, 0.5930157, 0.5943638, 
    0.5935606, 0.5906379, 0.6000335, 0.5951911, 0.6041679, 0.6015183, 
    0.6092895, 0.6054103, 0.6130582, 0.616364, 0.6194943, 0.6231793, 
    0.5928306, 0.5918136, 0.5936357, 0.5961673, 0.5985264, 0.6016796, 
    0.6020032, 0.6025964, 0.604136, 0.6054341, 0.6027843, 0.60576, 0.5946774, 
    0.6004559, 0.5914299, 0.5941321, 0.5960177, 0.5951895, 0.5995038, 
    0.6005259, 0.6047001, 0.6025379, 0.6155463, 0.60975, 0.6260031, 
    0.6214069, 0.5914588, 0.592827, 0.5976165, 0.5953323, 0.6018906, 
    0.6035177, 0.604844, 0.6065448, 0.6067286, 0.6077392, 0.6060841, 
    0.6076736, 0.6016863, 0.6043533, 0.5970665, 0.5988309, 0.5980185, 
    0.5971288, 0.5998793, 0.6028261, 0.6028888, 0.6038374, 0.6065205, 
    0.6019173, 0.6163, 0.6073706, 0.5943229, 0.596976, 0.5973556, 0.5963256, 
    0.6033544, 0.6007968, 0.6077145, 0.6058357, 0.6089177, 0.6073838, 
    0.6071586, 0.6051962, 0.6039783, 0.6009138, 0.5984336, 0.5964749, 
    0.5969296, 0.5990835, 0.6030067, 0.6067454, 0.6059241, 0.6086828, 
    0.6014124, 0.6044487, 0.6032732, 0.6063439, 0.5996386, 0.6053442, 
    0.5981902, 0.5988135, 0.6007462, 0.6046556, 0.6055239, 0.6064534, 
    0.6058796, 0.6031066, 0.6026536, 0.600699, 0.6001608, 0.5986778, 
    0.5974532, 0.598572, 0.5997495, 0.6031076, 0.6061528, 0.6094934, 
    0.6103142, 0.6142529, 0.6110448, 0.6163503, 0.6118369, 0.6196756, 
    0.6056762, 0.611704, 0.6008341, 0.6019941, 0.6040993, 0.6089594, 
    0.6063294, 0.6094063, 0.6026358, 0.5991582, 0.5982617, 0.5965938, 
    0.5982998, 0.5981609, 0.5997981, 0.5992714, 0.6032195, 0.601095, 
    0.6071531, 0.6093818, 0.6157289, 0.6196603, 0.6236942, 0.6254861, 
    0.6260328, 0.6262615,
  0.662225, 0.6677868, 0.6666974, 0.6712427, 0.6687127, 0.6717014, 0.6633441, 
    0.6680099, 0.665023, 0.6627212, 0.680266, 0.671447, 0.6897113, 0.683875, 
    0.6987641, 0.6887957, 0.7008164, 0.698471, 0.7055875, 0.7035305, 
    0.7128335, 0.706542, 0.7177785, 0.7113178, 0.712319, 0.7063369, 
    0.6732004, 0.6791539, 0.6728516, 0.6736922, 0.6733146, 0.6687649, 
    0.6664983, 0.6618037, 0.6626505, 0.6661009, 0.674071, 0.6713414, 
    0.6782679, 0.6781096, 0.6860121, 0.6824228, 0.6960331, 0.6920994, 
    0.703616, 0.700676, 0.7034774, 0.7026249, 0.7034885, 0.6991888, 
    0.7010232, 0.6972683, 0.6830918, 0.6871873, 0.6751373, 0.6681207, 
    0.6635474, 0.6603436, 0.6607946, 0.6616561, 0.6661212, 0.6703797, 
    0.673666, 0.6758847, 0.6780869, 0.6848563, 0.6885019, 0.6968353, 
    0.695313, 0.6978962, 0.7003852, 0.704614, 0.7039136, 0.7057922, 
    0.6978274, 0.7030962, 0.6944495, 0.6967888, 0.6786906, 0.6720753, 
    0.6693089, 0.6669066, 0.6611418, 0.6651112, 0.6635403, 0.6672907, 
    0.6696983, 0.668505, 0.6759456, 0.673031, 0.6887194, 0.6818594, 
    0.7000937, 0.6956248, 0.7011753, 0.6983294, 0.7032232, 0.6988151, 
    0.7064945, 0.7081947, 0.7070318, 0.7115247, 0.6985728, 0.7034776, 
    0.6684718, 0.6686661, 0.6695726, 0.6656078, 0.6653668, 0.6617806, 
    0.6649694, 0.6663377, 0.6698383, 0.6719286, 0.6739291, 0.6783752, 
    0.6834211, 0.6906249, 0.6959124, 0.6995118, 0.6972992, 0.6992517, 
    0.6970699, 0.696053, 0.7075566, 0.7010404, 0.7108741, 0.7103208, 
    0.7058372, 0.7103831, 0.6688025, 0.6676857, 0.6638407, 0.6668457, 
    0.6613926, 0.6644331, 0.6661955, 0.6730921, 0.6746283, 0.6760604, 
    0.6789089, 0.6826055, 0.6892046, 0.6950702, 0.7005305, 0.7001269, 
    0.700269, 0.7015022, 0.6984574, 0.7020051, 0.7026052, 0.7010394, 
    0.7102469, 0.7075857, 0.7103091, 0.7085731, 0.6680483, 0.6699319, 
    0.6689126, 0.6708323, 0.6694788, 0.6755452, 0.6773883, 0.6861677, 
    0.6825324, 0.6883389, 0.6831169, 0.6840355, 0.6885312, 0.6833965, 
    0.6947441, 0.6870037, 0.7015502, 0.6936396, 0.7020534, 0.7005067, 
    0.7030718, 0.7053891, 0.708331, 0.7138419, 0.7125561, 0.7172271, 
    0.6727619, 0.6752464, 0.6750264, 0.6776465, 0.6795993, 0.6838762, 
    0.690869, 0.6882196, 0.6931018, 0.694092, 0.6866816, 0.6912094, 
    0.6769204, 0.679183, 0.6778335, 0.6729574, 0.6888286, 0.6805772, 
    0.6960006, 0.6913904, 0.7050576, 0.6981798, 0.7118508, 0.7179043, 
    0.7237218, 0.7306814, 0.6766106, 0.6749126, 0.6779595, 0.6822281, 
    0.6862437, 0.6916696, 0.6922303, 0.6932602, 0.6959448, 0.6982216, 
    0.6935871, 0.6987951, 0.679711, 0.6895557, 0.6742734, 0.6787932, 
    0.6819746, 0.6805744, 0.6879182, 0.6896763, 0.6969326, 0.6931586, 
    0.7163985, 0.7058816, 0.7360994, 0.7273186, 0.6743217, 0.6766046, 
    0.6846904, 0.6808155, 0.6920352, 0.6948647, 0.697185, 0.7001794, 
    0.7005042, 0.7022953, 0.6993663, 0.7021788, 0.6916813, 0.6963251, 
    0.6837544, 0.6867647, 0.6853759, 0.6838603, 0.6885634, 0.6936595, 
    0.6937687, 0.6954227, 0.7001365, 0.6920815, 0.7177864, 0.701641, 
    0.6791142, 0.6836005, 0.6842462, 0.6824965, 0.6945798, 0.6901435, 
    0.7022514, 0.6989284, 0.7043933, 0.7016647, 0.7012655, 0.6978033, 
    0.6956689, 0.6903456, 0.6860849, 0.6827495, 0.6835217, 0.6871973, 
    0.693974, 0.700534, 0.6990843, 0.7039743, 0.6912071, 0.6964921, 
    0.6944382, 0.6998247, 0.6881497, 0.6980636, 0.6856692, 0.6867349, 
    0.6900561, 0.6968546, 0.6983795, 0.700018, 0.6990057, 0.694148, 
    0.6933596, 0.6899748, 0.6890475, 0.6865025, 0.6844124, 0.6863216, 
    0.6883402, 0.6941498, 0.6994875, 0.7054223, 0.7068934, 0.7140279, 
    0.7082076, 0.7178791, 0.709637, 0.7240613, 0.6986476, 0.7093968, 
    0.690208, 0.6922146, 0.6958805, 0.7044677, 0.6997991, 0.7052664, 
    0.6933287, 0.6873253, 0.6857911, 0.6829513, 0.6858563, 0.6856189, 
    0.6884237, 0.6875194, 0.6943446, 0.6906585, 0.7012556, 0.7052225, 
    0.7167342, 0.7240328, 0.7316638, 0.7351018, 0.7361567, 0.736599,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 XSMRPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 XSMRPOOL_RECOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZBOT =
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5 ;

 ZWT =
  8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882 ;

 ZWT_CH4_UNSAT =
  0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01893771, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01193812, 0.01893771, 
    0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01893771, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01893771, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01893771, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01193812, 0.01193812, 0.01193812, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01193812, 0.01193812, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01988501, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01193812, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 0.01988501, 
    0.01893771, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01893771, 
    0.01988501, 0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01893771, 
    0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01193812, 0.01893771, 0.01193812, 
    0.01893771, 0.01893771, 0.01988501, 0.01893771, 0.01893771, 0.01893771, 
    0.01893771, 0.01893771, 0.01893771, 0.01988501, 0.01988501, 0.01988501, 
    0.01988501, 0.01988501, 0.01988501, 0.01988501, 0.01893771, 0.01988501, 
    0.01893771, 0.01893771, 0.01893771, 0.01193812, 0.01193812, 0.01193812, 
    0.01193812, 0.01193812 ;

 ZWT_PERCH =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 o2_decomp_depth_unsat =
  3.353658e-11, 3.368474e-11, 3.365585e-11, 3.377543e-11, 3.370904e-11, 
    3.37873e-11, 3.356644e-11, 3.369039e-11, 3.36112e-11, 3.354962e-11, 
    3.400745e-11, 3.378049e-11, 3.424349e-11, 3.409845e-11, 3.446284e-11, 
    3.422082e-11, 3.451165e-11, 3.445576e-11, 3.462385e-11, 3.457562e-11, 
    3.479075e-11, 3.464599e-11, 3.490233e-11, 3.47561e-11, 3.477893e-11, 
    3.464105e-11, 3.382638e-11, 3.397943e-11, 3.381725e-11, 3.383907e-11, 
    3.382924e-11, 3.371027e-11, 3.365036e-11, 3.352495e-11, 3.354766e-11, 
    3.363974e-11, 3.384863e-11, 3.377762e-11, 3.395646e-11, 3.395243e-11, 
    3.415173e-11, 3.406181e-11, 3.439721e-11, 3.430176e-11, 3.457759e-11, 
    3.450812e-11, 3.457426e-11, 3.455414e-11, 3.457442e-11, 3.447263e-11, 
    3.451616e-11, 3.442662e-11, 3.407906e-11, 3.41813e-11, 3.387637e-11, 
    3.369325e-11, 3.357173e-11, 3.348559e-11, 3.349769e-11, 3.352092e-11, 
    3.364021e-11, 3.375245e-11, 3.383806e-11, 3.389531e-11, 3.395175e-11, 
    3.412284e-11, 3.421341e-11, 3.441643e-11, 3.437975e-11, 3.444182e-11, 
    3.450117e-11, 3.460084e-11, 3.458441e-11, 3.462831e-11, 3.444e-11, 
    3.45651e-11, 3.435858e-11, 3.441502e-11, 3.396745e-11, 3.379692e-11, 
    3.37245e-11, 3.366109e-11, 3.350703e-11, 3.361338e-11, 3.357141e-11, 
    3.367113e-11, 3.373455e-11, 3.370312e-11, 3.389684e-11, 3.382144e-11, 
    3.421873e-11, 3.404748e-11, 3.449429e-11, 3.43872e-11, 3.451986e-11, 
    3.445214e-11, 3.456813e-11, 3.446367e-11, 3.46446e-11, 3.468404e-11, 
    3.465701e-11, 3.476057e-11, 3.445767e-11, 3.457391e-11, 3.370244e-11, 
    3.370756e-11, 3.373136e-11, 3.362654e-11, 3.362012e-11, 3.352412e-11, 
    3.360945e-11, 3.364582e-11, 3.373813e-11, 3.379273e-11, 3.384466e-11, 
    3.3959e-11, 3.408673e-11, 3.426552e-11, 3.43941e-11, 3.44803e-11, 
    3.442739e-11, 3.447403e-11, 3.442182e-11, 3.43973e-11, 3.466916e-11, 
    3.451643e-11, 3.474557e-11, 3.473289e-11, 3.462908e-11, 3.473422e-11, 
    3.371109e-11, 3.368159e-11, 3.35794e-11, 3.36593e-11, 3.351361e-11, 
    3.359513e-11, 3.364197e-11, 3.382297e-11, 3.386273e-11, 3.389965e-11, 
    3.397255e-11, 3.406615e-11, 3.423056e-11, 3.437368e-11, 3.450449e-11, 
    3.449485e-11, 3.449821e-11, 3.452739e-11, 3.445496e-11, 3.453921e-11, 
    3.455332e-11, 3.451633e-11, 3.473109e-11, 3.466969e-11, 3.473248e-11, 
    3.469244e-11, 3.369112e-11, 3.374062e-11, 3.37138e-11, 3.376416e-11, 
    3.372861e-11, 3.388642e-11, 3.393372e-11, 3.415538e-11, 3.40643e-11, 
    3.420921e-11, 3.407895e-11, 3.410202e-11, 3.421382e-11, 3.408589e-11, 
    3.436568e-11, 3.417588e-11, 3.452849e-11, 3.433878e-11, 3.454031e-11, 
    3.450364e-11, 3.456423e-11, 3.461856e-11, 3.468684e-11, 3.481307e-11, 
    3.478375e-11, 3.488936e-11, 3.381447e-11, 3.387874e-11, 3.387306e-11, 
    3.394034e-11, 3.399011e-11, 3.409814e-11, 3.42715e-11, 3.420621e-11, 
    3.432594e-11, 3.435e-11, 3.416797e-11, 3.427967e-11, 3.392145e-11, 
    3.397921e-11, 3.394477e-11, 3.381902e-11, 3.422096e-11, 3.40145e-11, 
    3.439581e-11, 3.42838e-11, 3.461071e-11, 3.444803e-11, 3.476764e-11, 
    3.490448e-11, 3.503331e-11, 3.518397e-11, 3.391381e-11, 3.387004e-11, 
    3.394828e-11, 3.405666e-11, 3.415719e-11, 3.429105e-11, 3.43047e-11, 
    3.432974e-11, 3.439469e-11, 3.444937e-11, 3.433759e-11, 3.446298e-11, 
    3.399258e-11, 3.423888e-11, 3.385307e-11, 3.396915e-11, 3.404978e-11, 
    3.401438e-11, 3.419831e-11, 3.424165e-11, 3.441803e-11, 3.432683e-11, 
    3.48706e-11, 3.462978e-11, 3.529873e-11, 3.511154e-11, 3.385473e-11, 
    3.391352e-11, 3.41184e-11, 3.402087e-11, 3.429989e-11, 3.436865e-11, 
    3.44245e-11, 3.449602e-11, 3.450367e-11, 3.454606e-11, 3.447653e-11, 
    3.454325e-11, 3.429096e-11, 3.440362e-11, 3.409459e-11, 3.416969e-11, 
    3.41351e-11, 3.409712e-11, 3.421414e-11, 3.433896e-11, 3.434159e-11, 
    3.438156e-11, 3.449442e-11, 3.430038e-11, 3.490157e-11, 3.452998e-11, 
    3.397766e-11, 3.409104e-11, 3.41072e-11, 3.406325e-11, 3.436167e-11, 
    3.425346e-11, 3.454503e-11, 3.446611e-11, 3.45953e-11, 3.453108e-11, 
    3.452155e-11, 3.44391e-11, 3.438771e-11, 3.425815e-11, 3.415271e-11, 
    3.406922e-11, 3.408855e-11, 3.41803e-11, 3.43465e-11, 3.450394e-11, 
    3.446939e-11, 3.458504e-11, 3.427893e-11, 3.44072e-11, 3.435755e-11, 
    3.448688e-11, 3.420434e-11, 3.444553e-11, 3.414271e-11, 3.416918e-11, 
    3.425121e-11, 3.441643e-11, 3.445293e-11, 3.4492e-11, 3.446782e-11, 
    3.435098e-11, 3.43318e-11, 3.424899e-11, 3.42261e-11, 3.41631e-11, 
    3.411086e-11, 3.415852e-11, 3.42085e-11, 3.435075e-11, 3.447898e-11, 
    3.46189e-11, 3.465316e-11, 3.481683e-11, 3.468353e-11, 3.490347e-11, 
    3.47164e-11, 3.504027e-11, 3.445941e-11, 3.471161e-11, 3.425496e-11, 
    3.430404e-11, 3.439291e-11, 3.459695e-11, 3.448669e-11, 3.46156e-11, 
    3.433102e-11, 3.418352e-11, 3.414535e-11, 3.407425e-11, 3.414691e-11, 
    3.4141e-11, 3.421059e-11, 3.418815e-11, 3.435538e-11, 3.426551e-11, 
    3.452085e-11, 3.461417e-11, 3.487789e-11, 3.503972e-11, 3.520463e-11, 
    3.527744e-11, 3.52996e-11, 3.530884e-11,
  1.907281e-11, 1.921687e-11, 1.918884e-11, 1.930526e-11, 1.924065e-11, 
    1.931692e-11, 1.910199e-11, 1.92226e-11, 1.914557e-11, 1.908577e-11, 
    1.953193e-11, 1.931046e-11, 1.976297e-11, 1.9621e-11, 1.997833e-11, 
    1.974085e-11, 2.002633e-11, 1.997147e-11, 2.013679e-11, 2.008938e-11, 
    2.030135e-11, 2.015868e-11, 2.041155e-11, 2.026725e-11, 2.02898e-11, 
    2.015398e-11, 1.935496e-11, 1.95043e-11, 1.934612e-11, 1.936739e-11, 
    1.935785e-11, 1.924198e-11, 1.918368e-11, 1.906182e-11, 1.908392e-11, 
    1.917344e-11, 1.937695e-11, 1.930778e-11, 1.948229e-11, 1.947835e-11, 
    1.967328e-11, 1.95853e-11, 1.9914e-11, 1.982038e-11, 2.009135e-11, 
    2.002308e-11, 2.008814e-11, 2.006841e-11, 2.00884e-11, 1.99883e-11, 
    2.003117e-11, 1.994317e-11, 1.960177e-11, 1.970188e-11, 1.940384e-11, 
    1.922543e-11, 1.910727e-11, 1.902359e-11, 1.903541e-11, 1.905795e-11, 
    1.917396e-11, 1.928328e-11, 1.936674e-11, 1.942264e-11, 1.947778e-11, 
    1.964501e-11, 1.973375e-11, 1.993295e-11, 1.989695e-11, 1.995795e-11, 
    2.001629e-11, 2.011438e-11, 2.009823e-11, 2.014148e-11, 1.995634e-11, 
    2.007932e-11, 1.987646e-11, 1.993186e-11, 1.949276e-11, 1.932644e-11, 
    1.925589e-11, 1.919422e-11, 1.90445e-11, 1.914785e-11, 1.910708e-11, 
    1.920412e-11, 1.926588e-11, 1.923533e-11, 1.942417e-11, 1.935067e-11, 
    1.973901e-11, 1.95714e-11, 2.000949e-11, 1.990433e-11, 2.003472e-11, 
    1.996815e-11, 2.008226e-11, 1.997955e-11, 2.015759e-11, 2.019643e-11, 
    2.016989e-11, 2.027193e-11, 1.997386e-11, 2.008814e-11, 1.923447e-11, 
    1.923945e-11, 1.926267e-11, 1.91607e-11, 1.915447e-11, 1.906121e-11, 
    1.914418e-11, 1.917955e-11, 1.926946e-11, 1.932271e-11, 1.937338e-11, 
    1.948496e-11, 1.960985e-11, 1.978498e-11, 1.991114e-11, 1.999588e-11, 
    1.994391e-11, 1.998979e-11, 1.99385e-11, 1.991448e-11, 2.018187e-11, 
    2.003157e-11, 2.025724e-11, 2.024473e-11, 2.014251e-11, 2.024614e-11, 
    1.924295e-11, 1.921429e-11, 1.91149e-11, 1.919266e-11, 1.905107e-11, 
    1.913028e-11, 1.917587e-11, 1.93522e-11, 1.939103e-11, 1.942705e-11, 
    1.949827e-11, 1.95898e-11, 1.975075e-11, 1.989118e-11, 2.001969e-11, 
    2.001026e-11, 2.001358e-11, 2.004233e-11, 1.997115e-11, 2.005402e-11, 
    2.006794e-11, 2.003155e-11, 2.024306e-11, 2.018255e-11, 2.024447e-11, 
    2.020506e-11, 1.92236e-11, 1.927185e-11, 1.924577e-11, 1.929482e-11, 
    1.926026e-11, 1.941409e-11, 1.94603e-11, 1.967706e-11, 1.9588e-11, 
    1.972981e-11, 1.960239e-11, 1.962494e-11, 1.973444e-11, 1.960927e-11, 
    1.988342e-11, 1.96974e-11, 2.004344e-11, 1.985713e-11, 2.005514e-11, 
    2.001913e-11, 2.007876e-11, 2.013222e-11, 2.019955e-11, 2.032398e-11, 
    2.029514e-11, 2.039936e-11, 1.934385e-11, 1.940658e-11, 1.940106e-11, 
    1.946678e-11, 1.951543e-11, 1.962104e-11, 1.979086e-11, 1.972694e-11, 
    1.984434e-11, 1.986794e-11, 1.96896e-11, 1.979903e-11, 1.944861e-11, 
    1.950506e-11, 1.947145e-11, 1.93488e-11, 1.974166e-11, 1.953968e-11, 
    1.991323e-11, 1.980338e-11, 2.01246e-11, 1.996461e-11, 2.027927e-11, 
    2.041432e-11, 2.054171e-11, 2.069093e-11, 1.944085e-11, 1.939819e-11, 
    1.94746e-11, 1.958049e-11, 1.967893e-11, 1.981008e-11, 1.982351e-11, 
    1.984812e-11, 1.991192e-11, 1.996561e-11, 1.98559e-11, 1.997908e-11, 
    1.951816e-11, 1.975923e-11, 1.938207e-11, 1.949536e-11, 1.957424e-11, 
    1.953963e-11, 1.971964e-11, 1.976215e-11, 1.993524e-11, 1.98457e-11, 
    2.038095e-11, 2.014351e-11, 2.08048e-11, 2.061925e-11, 1.93833e-11, 
    1.944071e-11, 1.964099e-11, 1.95456e-11, 1.981884e-11, 1.98863e-11, 
    1.994122e-11, 2.001148e-11, 2.001907e-11, 2.006076e-11, 1.999247e-11, 
    2.005806e-11, 1.981035e-11, 1.992091e-11, 1.961806e-11, 1.969161e-11, 
    1.965776e-11, 1.962066e-11, 1.973526e-11, 1.985763e-11, 1.986025e-11, 
    1.989954e-11, 2.001041e-11, 1.981995e-11, 2.041166e-11, 2.004549e-11, 
    1.950338e-11, 1.961425e-11, 1.963011e-11, 1.958712e-11, 1.987954e-11, 
    1.977341e-11, 2.005974e-11, 1.998221e-11, 2.01093e-11, 2.004611e-11, 
    2.003682e-11, 1.995578e-11, 1.990538e-11, 1.977827e-11, 1.967506e-11, 
    1.959336e-11, 1.961234e-11, 1.970213e-11, 1.986512e-11, 2.001976e-11, 
    1.998585e-11, 2.009963e-11, 1.979898e-11, 1.992485e-11, 1.987617e-11, 
    2.00032e-11, 1.972524e-11, 1.996183e-11, 1.966493e-11, 1.969089e-11, 
    1.97713e-11, 1.993339e-11, 1.996932e-11, 2.000771e-11, 1.998402e-11, 
    1.986927e-11, 1.985049e-11, 1.976935e-11, 1.974696e-11, 1.968524e-11, 
    1.963419e-11, 1.968083e-11, 1.972985e-11, 1.986932e-11, 1.99953e-11, 
    2.013298e-11, 2.016673e-11, 2.032811e-11, 2.01967e-11, 2.041371e-11, 
    2.022914e-11, 2.054901e-11, 1.997558e-11, 2.022374e-11, 1.977496e-11, 
    1.982314e-11, 1.991037e-11, 2.011099e-11, 2.00026e-11, 2.012938e-11, 
    1.984976e-11, 1.970523e-11, 1.96679e-11, 1.959832e-11, 1.966949e-11, 
    1.96637e-11, 1.973188e-11, 1.970996e-11, 1.987395e-11, 1.97858e-11, 
    2.003658e-11, 2.012838e-11, 2.038843e-11, 2.054843e-11, 2.071176e-11, 
    2.0784e-11, 2.080601e-11, 2.081521e-11,
  1.783539e-11, 1.799306e-11, 1.796236e-11, 1.808986e-11, 1.801909e-11, 
    1.810264e-11, 1.786731e-11, 1.799933e-11, 1.791501e-11, 1.784957e-11, 
    1.833837e-11, 1.809556e-11, 1.859205e-11, 1.843613e-11, 1.882885e-11, 
    1.856774e-11, 1.888168e-11, 1.88213e-11, 1.90033e-11, 1.895109e-11, 
    1.918465e-11, 1.902742e-11, 1.93062e-11, 1.914705e-11, 1.917191e-11, 
    1.902224e-11, 1.814432e-11, 1.830806e-11, 1.813463e-11, 1.815794e-11, 
    1.814748e-11, 1.802055e-11, 1.795672e-11, 1.782337e-11, 1.784755e-11, 
    1.794551e-11, 1.816843e-11, 1.809263e-11, 1.828392e-11, 1.827959e-11, 
    1.849353e-11, 1.839694e-11, 1.875808e-11, 1.865514e-11, 1.895326e-11, 
    1.88781e-11, 1.894973e-11, 1.8928e-11, 1.895001e-11, 1.883983e-11, 
    1.8887e-11, 1.879017e-11, 1.841501e-11, 1.852494e-11, 1.81979e-11, 
    1.800242e-11, 1.787309e-11, 1.778156e-11, 1.779449e-11, 1.781914e-11, 
    1.794608e-11, 1.806578e-11, 1.815723e-11, 1.821851e-11, 1.827897e-11, 
    1.846249e-11, 1.855995e-11, 1.877892e-11, 1.873933e-11, 1.880643e-11, 
    1.887063e-11, 1.897862e-11, 1.896083e-11, 1.900847e-11, 1.880466e-11, 
    1.894001e-11, 1.871679e-11, 1.877773e-11, 1.829541e-11, 1.811306e-11, 
    1.803578e-11, 1.796826e-11, 1.780443e-11, 1.79175e-11, 1.787289e-11, 
    1.79791e-11, 1.804672e-11, 1.801326e-11, 1.822018e-11, 1.813962e-11, 
    1.856573e-11, 1.838168e-11, 1.886314e-11, 1.874745e-11, 1.889091e-11, 
    1.881765e-11, 1.894325e-11, 1.88302e-11, 1.902621e-11, 1.9069e-11, 
    1.903976e-11, 1.915221e-11, 1.882394e-11, 1.894973e-11, 1.801233e-11, 
    1.801778e-11, 1.80432e-11, 1.793156e-11, 1.792474e-11, 1.782271e-11, 
    1.791349e-11, 1.79522e-11, 1.805065e-11, 1.810898e-11, 1.816451e-11, 
    1.828685e-11, 1.842389e-11, 1.861624e-11, 1.875494e-11, 1.884816e-11, 
    1.879098e-11, 1.884146e-11, 1.878503e-11, 1.875861e-11, 1.905296e-11, 
    1.888744e-11, 1.913602e-11, 1.912223e-11, 1.90096e-11, 1.912379e-11, 
    1.802161e-11, 1.799023e-11, 1.788144e-11, 1.796655e-11, 1.781161e-11, 
    1.789827e-11, 1.794817e-11, 1.81413e-11, 1.818385e-11, 1.822334e-11, 
    1.830144e-11, 1.840188e-11, 1.857863e-11, 1.873299e-11, 1.887437e-11, 
    1.8864e-11, 1.886765e-11, 1.889929e-11, 1.882096e-11, 1.891216e-11, 
    1.892748e-11, 1.888743e-11, 1.912038e-11, 1.905371e-11, 1.912194e-11, 
    1.907851e-11, 1.800043e-11, 1.805326e-11, 1.80247e-11, 1.807842e-11, 
    1.804057e-11, 1.820913e-11, 1.82598e-11, 1.849768e-11, 1.83999e-11, 
    1.855562e-11, 1.841569e-11, 1.844045e-11, 1.85607e-11, 1.842325e-11, 
    1.872446e-11, 1.852002e-11, 1.890052e-11, 1.869555e-11, 1.891339e-11, 
    1.887376e-11, 1.89394e-11, 1.899827e-11, 1.907244e-11, 1.92096e-11, 
    1.91778e-11, 1.929275e-11, 1.813215e-11, 1.82009e-11, 1.819485e-11, 
    1.826691e-11, 1.832027e-11, 1.843617e-11, 1.86227e-11, 1.855246e-11, 
    1.868149e-11, 1.870743e-11, 1.851145e-11, 1.863168e-11, 1.824698e-11, 
    1.83089e-11, 1.827202e-11, 1.813757e-11, 1.856863e-11, 1.834688e-11, 
    1.875724e-11, 1.863646e-11, 1.898987e-11, 1.881376e-11, 1.916031e-11, 
    1.930925e-11, 1.944987e-11, 1.961472e-11, 1.823847e-11, 1.819171e-11, 
    1.827548e-11, 1.839165e-11, 1.849973e-11, 1.864382e-11, 1.865859e-11, 
    1.868564e-11, 1.875579e-11, 1.881486e-11, 1.86942e-11, 1.882968e-11, 
    1.832327e-11, 1.858794e-11, 1.817403e-11, 1.829825e-11, 1.83848e-11, 
    1.834682e-11, 1.854444e-11, 1.859115e-11, 1.878145e-11, 1.868298e-11, 
    1.927244e-11, 1.901071e-11, 1.974063e-11, 1.953551e-11, 1.817538e-11, 
    1.823831e-11, 1.845806e-11, 1.835337e-11, 1.865345e-11, 1.872763e-11, 
    1.878802e-11, 1.886534e-11, 1.887369e-11, 1.891957e-11, 1.884441e-11, 
    1.89166e-11, 1.864412e-11, 1.876569e-11, 1.84329e-11, 1.851366e-11, 
    1.847649e-11, 1.843575e-11, 1.856161e-11, 1.869609e-11, 1.869897e-11, 
    1.874218e-11, 1.886416e-11, 1.865467e-11, 1.930632e-11, 1.890277e-11, 
    1.830705e-11, 1.842872e-11, 1.844613e-11, 1.839894e-11, 1.872019e-11, 
    1.860352e-11, 1.891846e-11, 1.883312e-11, 1.897302e-11, 1.890345e-11, 
    1.889322e-11, 1.880404e-11, 1.874861e-11, 1.860886e-11, 1.849548e-11, 
    1.840578e-11, 1.842662e-11, 1.852521e-11, 1.870433e-11, 1.887445e-11, 
    1.883713e-11, 1.896238e-11, 1.863163e-11, 1.877002e-11, 1.871648e-11, 
    1.885622e-11, 1.85506e-11, 1.88107e-11, 1.848435e-11, 1.851287e-11, 
    1.860121e-11, 1.877942e-11, 1.881895e-11, 1.886119e-11, 1.883512e-11, 
    1.870889e-11, 1.868825e-11, 1.859906e-11, 1.857446e-11, 1.850666e-11, 
    1.845061e-11, 1.850182e-11, 1.855566e-11, 1.870894e-11, 1.884753e-11, 
    1.899911e-11, 1.903628e-11, 1.921415e-11, 1.90693e-11, 1.930857e-11, 
    1.910505e-11, 1.945793e-11, 1.882583e-11, 1.909909e-11, 1.860523e-11, 
    1.865818e-11, 1.87541e-11, 1.897488e-11, 1.885556e-11, 1.899514e-11, 
    1.868744e-11, 1.852861e-11, 1.848762e-11, 1.841123e-11, 1.848937e-11, 
    1.848301e-11, 1.85579e-11, 1.853382e-11, 1.871404e-11, 1.861714e-11, 
    1.889296e-11, 1.899404e-11, 1.928069e-11, 1.945728e-11, 1.963774e-11, 
    1.971762e-11, 1.974196e-11, 1.975214e-11,
  1.829493e-11, 1.846855e-11, 1.843474e-11, 1.857523e-11, 1.849723e-11, 
    1.858931e-11, 1.833006e-11, 1.847546e-11, 1.838258e-11, 1.831052e-11, 
    1.884933e-11, 1.858151e-11, 1.912946e-11, 1.895722e-11, 1.939129e-11, 
    1.910261e-11, 1.944975e-11, 1.938293e-11, 1.958437e-11, 1.952656e-11, 
    1.97853e-11, 1.961108e-11, 1.992006e-11, 1.974363e-11, 1.977118e-11, 
    1.960535e-11, 1.863525e-11, 1.881588e-11, 1.862458e-11, 1.865028e-11, 
    1.863874e-11, 1.849884e-11, 1.842853e-11, 1.828169e-11, 1.830831e-11, 
    1.841618e-11, 1.866184e-11, 1.857827e-11, 1.878922e-11, 1.878445e-11, 
    1.902061e-11, 1.891396e-11, 1.9313e-11, 1.919918e-11, 1.952897e-11, 
    1.944578e-11, 1.952506e-11, 1.9501e-11, 1.952537e-11, 1.940343e-11, 
    1.945564e-11, 1.93485e-11, 1.893391e-11, 1.905531e-11, 1.869434e-11, 
    1.847888e-11, 1.833643e-11, 1.823567e-11, 1.82499e-11, 1.827704e-11, 
    1.841681e-11, 1.854869e-11, 1.864949e-11, 1.871706e-11, 1.878376e-11, 
    1.898635e-11, 1.909399e-11, 1.933606e-11, 1.929226e-11, 1.936648e-11, 
    1.943751e-11, 1.955705e-11, 1.953735e-11, 1.95901e-11, 1.936452e-11, 
    1.95143e-11, 1.926734e-11, 1.933474e-11, 1.880192e-11, 1.86008e-11, 
    1.851563e-11, 1.844123e-11, 1.826084e-11, 1.838533e-11, 1.833621e-11, 
    1.845317e-11, 1.852768e-11, 1.849081e-11, 1.871891e-11, 1.863007e-11, 
    1.910037e-11, 1.889711e-11, 1.942922e-11, 1.930125e-11, 1.945996e-11, 
    1.937889e-11, 1.951789e-11, 1.939277e-11, 1.960975e-11, 1.965715e-11, 
    1.962475e-11, 1.974934e-11, 1.938585e-11, 1.952506e-11, 1.848978e-11, 
    1.849579e-11, 1.85238e-11, 1.840081e-11, 1.83933e-11, 1.828096e-11, 
    1.838091e-11, 1.842355e-11, 1.8532e-11, 1.85963e-11, 1.865752e-11, 
    1.879246e-11, 1.894371e-11, 1.915619e-11, 1.930953e-11, 1.941265e-11, 
    1.934939e-11, 1.940523e-11, 1.934281e-11, 1.931358e-11, 1.963938e-11, 
    1.945612e-11, 1.97314e-11, 1.971611e-11, 1.959135e-11, 1.971784e-11, 
    1.850001e-11, 1.846543e-11, 1.834562e-11, 1.843935e-11, 1.826875e-11, 
    1.836415e-11, 1.841911e-11, 1.863193e-11, 1.867884e-11, 1.87224e-11, 
    1.880856e-11, 1.891941e-11, 1.911462e-11, 1.928525e-11, 1.944165e-11, 
    1.943017e-11, 1.943421e-11, 1.946923e-11, 1.938255e-11, 1.948347e-11, 
    1.950044e-11, 1.94561e-11, 1.971407e-11, 1.96402e-11, 1.971579e-11, 
    1.966768e-11, 1.847667e-11, 1.853488e-11, 1.850342e-11, 1.856261e-11, 
    1.85209e-11, 1.870673e-11, 1.876262e-11, 1.90252e-11, 1.891722e-11, 
    1.90892e-11, 1.893466e-11, 1.8962e-11, 1.909483e-11, 1.894299e-11, 
    1.927583e-11, 1.904988e-11, 1.947059e-11, 1.924387e-11, 1.948484e-11, 
    1.944097e-11, 1.951362e-11, 1.95788e-11, 1.966095e-11, 1.981295e-11, 
    1.97777e-11, 1.990514e-11, 1.862184e-11, 1.869765e-11, 1.869097e-11, 
    1.877045e-11, 1.882934e-11, 1.895727e-11, 1.916332e-11, 1.908571e-11, 
    1.92283e-11, 1.925699e-11, 1.90404e-11, 1.917325e-11, 1.874847e-11, 
    1.881679e-11, 1.87761e-11, 1.862781e-11, 1.910358e-11, 1.88587e-11, 
    1.931207e-11, 1.917853e-11, 1.95695e-11, 1.93746e-11, 1.975831e-11, 
    1.992345e-11, 2.007945e-11, 2.026251e-11, 1.873909e-11, 1.86875e-11, 
    1.877991e-11, 1.890813e-11, 1.902746e-11, 1.918666e-11, 1.920299e-11, 
    1.92329e-11, 1.931047e-11, 1.937581e-11, 1.924236e-11, 1.93922e-11, 
    1.883266e-11, 1.912491e-11, 1.866802e-11, 1.880505e-11, 1.890056e-11, 
    1.885863e-11, 1.907685e-11, 1.912846e-11, 1.933886e-11, 1.922995e-11, 
    1.988263e-11, 1.959259e-11, 2.040242e-11, 2.017453e-11, 1.86695e-11, 
    1.873891e-11, 1.898145e-11, 1.886586e-11, 1.919731e-11, 1.927932e-11, 
    1.934611e-11, 1.943166e-11, 1.94409e-11, 1.949168e-11, 1.94085e-11, 
    1.948839e-11, 1.9187e-11, 1.932141e-11, 1.895365e-11, 1.904285e-11, 
    1.900179e-11, 1.89568e-11, 1.909581e-11, 1.924446e-11, 1.924764e-11, 
    1.929542e-11, 1.943038e-11, 1.919866e-11, 1.992022e-11, 1.947311e-11, 
    1.881474e-11, 1.894905e-11, 1.896826e-11, 1.891616e-11, 1.92711e-11, 
    1.914212e-11, 1.949044e-11, 1.939601e-11, 1.955085e-11, 1.947383e-11, 
    1.946251e-11, 1.936384e-11, 1.930252e-11, 1.914803e-11, 1.902276e-11, 
    1.892371e-11, 1.894672e-11, 1.90556e-11, 1.925357e-11, 1.944174e-11, 
    1.940044e-11, 1.953906e-11, 1.917319e-11, 1.93262e-11, 1.9267e-11, 
    1.942156e-11, 1.908365e-11, 1.937123e-11, 1.901047e-11, 1.904197e-11, 
    1.913957e-11, 1.933661e-11, 1.938032e-11, 1.942706e-11, 1.939822e-11, 
    1.925861e-11, 1.923578e-11, 1.913719e-11, 1.911002e-11, 1.903511e-11, 
    1.89732e-11, 1.902976e-11, 1.908925e-11, 1.925866e-11, 1.941195e-11, 
    1.957973e-11, 1.96209e-11, 1.981801e-11, 1.965748e-11, 1.992272e-11, 
    1.969712e-11, 2.008843e-11, 1.938795e-11, 1.96905e-11, 1.914401e-11, 
    1.920253e-11, 1.93086e-11, 1.955292e-11, 1.942083e-11, 1.957535e-11, 
    1.923488e-11, 1.905937e-11, 1.901408e-11, 1.892973e-11, 1.901601e-11, 
    1.900899e-11, 1.909171e-11, 1.906511e-11, 1.92643e-11, 1.915718e-11, 
    1.946223e-11, 1.957412e-11, 1.989177e-11, 2.00877e-11, 2.028808e-11, 
    2.037684e-11, 2.04039e-11, 2.041521e-11,
  1.973493e-11, 1.991887e-11, 1.988303e-11, 2.003195e-11, 1.994926e-11, 
    2.004689e-11, 1.977214e-11, 1.99262e-11, 1.982776e-11, 1.975144e-11, 
    2.032279e-11, 2.003861e-11, 2.062036e-11, 2.043734e-11, 2.089887e-11, 
    2.059183e-11, 2.096109e-11, 2.088996e-11, 2.110444e-11, 2.104287e-11, 
    2.131862e-11, 2.11329e-11, 2.146236e-11, 2.127417e-11, 2.130355e-11, 
    2.112679e-11, 2.00956e-11, 2.028729e-11, 2.008428e-11, 2.011154e-11, 
    2.009931e-11, 1.995097e-11, 1.987647e-11, 1.97209e-11, 1.974909e-11, 
    1.986337e-11, 2.012381e-11, 2.003517e-11, 2.025896e-11, 2.025389e-11, 
    2.050468e-11, 2.039138e-11, 2.081555e-11, 2.069448e-11, 2.104543e-11, 
    2.095685e-11, 2.104127e-11, 2.101565e-11, 2.10416e-11, 2.091178e-11, 
    2.096735e-11, 2.085331e-11, 2.041258e-11, 2.054155e-11, 2.015828e-11, 
    1.992983e-11, 1.977888e-11, 1.967217e-11, 1.968724e-11, 1.971598e-11, 
    1.986404e-11, 2.00038e-11, 2.01107e-11, 2.018239e-11, 2.025316e-11, 
    2.046829e-11, 2.058266e-11, 2.084008e-11, 2.079348e-11, 2.087246e-11, 
    2.094805e-11, 2.107534e-11, 2.105436e-11, 2.111055e-11, 2.087036e-11, 
    2.102982e-11, 2.076696e-11, 2.083867e-11, 2.027247e-11, 2.005906e-11, 
    1.996878e-11, 1.988992e-11, 1.969883e-11, 1.983068e-11, 1.977864e-11, 
    1.990256e-11, 1.998154e-11, 1.994245e-11, 2.018435e-11, 2.009011e-11, 
    2.058945e-11, 2.03735e-11, 2.093923e-11, 2.080304e-11, 2.097194e-11, 
    2.088565e-11, 2.103364e-11, 2.090043e-11, 2.113148e-11, 2.1182e-11, 
    2.114747e-11, 2.128025e-11, 2.089306e-11, 2.104127e-11, 1.994136e-11, 
    1.994773e-11, 1.997742e-11, 1.984709e-11, 1.983913e-11, 1.972013e-11, 
    1.982599e-11, 1.987117e-11, 1.998612e-11, 2.005429e-11, 2.011922e-11, 
    2.026239e-11, 2.042299e-11, 2.064877e-11, 2.081185e-11, 2.092158e-11, 
    2.085426e-11, 2.091369e-11, 2.084726e-11, 2.081616e-11, 2.116306e-11, 
    2.096787e-11, 2.126113e-11, 2.124484e-11, 2.111189e-11, 2.124667e-11, 
    1.99522e-11, 1.991555e-11, 1.978861e-11, 1.988791e-11, 1.97072e-11, 
    1.980824e-11, 1.986648e-11, 2.009209e-11, 2.014184e-11, 2.018805e-11, 
    2.027948e-11, 2.039717e-11, 2.060459e-11, 2.078603e-11, 2.095245e-11, 
    2.094023e-11, 2.094453e-11, 2.098182e-11, 2.088955e-11, 2.099699e-11, 
    2.101505e-11, 2.096784e-11, 2.124266e-11, 2.116393e-11, 2.124449e-11, 
    2.119321e-11, 1.992746e-11, 1.998917e-11, 1.995581e-11, 2.001858e-11, 
    1.997435e-11, 2.017144e-11, 2.023074e-11, 2.050956e-11, 2.039486e-11, 
    2.057757e-11, 2.041337e-11, 2.044241e-11, 2.058357e-11, 2.042222e-11, 
    2.077601e-11, 2.053579e-11, 2.098327e-11, 2.074202e-11, 2.099844e-11, 
    2.095173e-11, 2.102909e-11, 2.109852e-11, 2.118604e-11, 2.13481e-11, 
    2.13105e-11, 2.144643e-11, 2.008137e-11, 2.01618e-11, 2.01547e-11, 
    2.023904e-11, 2.030154e-11, 2.043738e-11, 2.065635e-11, 2.057385e-11, 
    2.072545e-11, 2.075596e-11, 2.05257e-11, 2.066691e-11, 2.021572e-11, 
    2.028823e-11, 2.024503e-11, 2.008772e-11, 2.059286e-11, 2.033272e-11, 
    2.081455e-11, 2.067252e-11, 2.108861e-11, 2.088109e-11, 2.128983e-11, 
    2.146598e-11, 2.16325e-11, 2.18281e-11, 2.020576e-11, 2.015102e-11, 
    2.024908e-11, 2.03852e-11, 2.051195e-11, 2.068117e-11, 2.069852e-11, 
    2.073033e-11, 2.081285e-11, 2.088237e-11, 2.074041e-11, 2.089982e-11, 
    2.030509e-11, 2.061552e-11, 2.013036e-11, 2.027577e-11, 2.037716e-11, 
    2.033264e-11, 2.056443e-11, 2.061928e-11, 2.084306e-11, 2.07272e-11, 
    2.142244e-11, 2.111321e-11, 2.197769e-11, 2.173408e-11, 2.013192e-11, 
    2.020556e-11, 2.046308e-11, 2.034032e-11, 2.069249e-11, 2.077972e-11, 
    2.085077e-11, 2.094182e-11, 2.095166e-11, 2.100572e-11, 2.091717e-11, 
    2.100222e-11, 2.068153e-11, 2.082449e-11, 2.043354e-11, 2.05283e-11, 
    2.048467e-11, 2.043688e-11, 2.058459e-11, 2.074264e-11, 2.074601e-11, 
    2.079684e-11, 2.09405e-11, 2.069392e-11, 2.146257e-11, 2.098599e-11, 
    2.028604e-11, 2.042866e-11, 2.044906e-11, 2.039372e-11, 2.077096e-11, 
    2.063382e-11, 2.10044e-11, 2.090387e-11, 2.106874e-11, 2.098672e-11, 
    2.097467e-11, 2.086963e-11, 2.080439e-11, 2.06401e-11, 2.050696e-11, 
    2.040174e-11, 2.042618e-11, 2.054186e-11, 2.075233e-11, 2.095256e-11, 
    2.09086e-11, 2.105618e-11, 2.066684e-11, 2.082959e-11, 2.076661e-11, 
    2.093107e-11, 2.057166e-11, 2.087754e-11, 2.04939e-11, 2.052737e-11, 
    2.06311e-11, 2.084067e-11, 2.088718e-11, 2.093693e-11, 2.090622e-11, 
    2.075768e-11, 2.07334e-11, 2.062857e-11, 2.059969e-11, 2.052008e-11, 
    2.045431e-11, 2.05144e-11, 2.057762e-11, 2.075774e-11, 2.092084e-11, 
    2.109951e-11, 2.114336e-11, 2.135351e-11, 2.118237e-11, 2.146524e-11, 
    2.122464e-11, 2.164212e-11, 2.089532e-11, 2.121756e-11, 2.063582e-11, 
    2.069804e-11, 2.081087e-11, 2.107096e-11, 2.09303e-11, 2.109484e-11, 
    2.073245e-11, 2.054587e-11, 2.049773e-11, 2.040813e-11, 2.049978e-11, 
    2.049232e-11, 2.058023e-11, 2.055195e-11, 2.076373e-11, 2.064982e-11, 
    2.097437e-11, 2.109354e-11, 2.143217e-11, 2.164132e-11, 2.185541e-11, 
    2.195033e-11, 2.197926e-11, 2.199137e-11,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
